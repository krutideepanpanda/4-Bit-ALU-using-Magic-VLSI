magic
tech scmos
timestamp 1636190380
<< ab >>
rect -271 85 -23 93
rect -271 59 -191 85
rect -265 55 -191 59
rect -271 53 -191 55
rect -190 53 -87 85
rect -86 53 -23 85
rect -271 21 -23 53
rect 5 56 55 105
rect 5 54 14 56
rect 16 54 34 56
rect 36 54 44 56
rect 46 54 55 56
rect 5 53 55 54
rect 105 56 155 105
rect 105 54 114 56
rect 116 54 134 56
rect 136 54 144 56
rect 146 54 155 56
rect -196 16 -190 21
rect -92 16 -86 21
rect 5 17 51 53
rect 5 5 55 17
rect 105 5 155 54
rect 201 5 321 105
<< nwell >>
rect -276 53 326 110
<< pwell >>
rect -276 0 326 53
<< poly >>
rect 40 99 42 103
rect 16 91 18 95
rect -249 87 -247 91
rect -242 87 -240 91
rect -262 77 -260 82
rect -174 87 -172 91
rect -222 78 -220 82
rect -212 80 -210 85
rect -202 80 -200 85
rect -262 56 -260 59
rect -249 56 -247 66
rect -242 63 -240 66
rect -242 61 -236 63
rect -242 59 -240 61
rect -238 59 -236 61
rect -242 57 -236 59
rect -262 54 -256 56
rect -262 52 -260 54
rect -258 52 -256 54
rect -262 50 -256 52
rect -252 54 -246 56
rect -252 52 -250 54
rect -248 52 -246 54
rect -252 50 -246 52
rect -262 47 -260 50
rect -252 47 -250 50
rect -242 47 -240 57
rect -222 56 -220 60
rect -212 56 -210 67
rect -202 64 -200 67
rect -202 62 -196 64
rect -202 60 -200 62
rect -198 60 -196 62
rect -202 58 -196 60
rect -189 62 -183 64
rect -189 60 -187 62
rect -185 60 -183 62
rect -138 87 -136 91
rect -158 78 -156 82
rect -148 78 -146 82
rect -70 87 -68 91
rect -118 78 -116 82
rect -108 80 -106 85
rect -98 80 -96 85
rect -189 58 -183 60
rect -222 54 -216 56
rect -222 52 -220 54
rect -218 52 -216 54
rect -222 50 -216 52
rect -212 54 -206 56
rect -212 52 -210 54
rect -208 52 -206 54
rect -212 50 -206 52
rect -222 45 -220 50
rect -209 45 -207 50
rect -202 45 -200 58
rect -185 57 -183 58
rect -174 57 -172 60
rect -158 57 -156 60
rect -185 55 -172 57
rect -166 55 -156 57
rect -148 56 -146 60
rect -138 57 -136 60
rect -182 47 -180 55
rect -166 51 -164 55
rect -173 49 -164 51
rect -152 54 -146 56
rect -152 52 -150 54
rect -148 52 -146 54
rect -152 50 -146 52
rect -142 55 -136 57
rect -142 53 -140 55
rect -138 53 -136 55
rect -142 51 -136 53
rect -118 56 -116 60
rect -108 56 -106 67
rect -98 64 -96 67
rect -98 62 -92 64
rect -98 60 -96 62
rect -94 60 -92 62
rect -98 58 -92 60
rect -85 62 -79 64
rect -85 60 -83 62
rect -81 60 -79 62
rect -34 87 -32 91
rect -54 78 -52 82
rect -44 78 -42 82
rect 28 90 30 94
rect 16 68 18 71
rect 12 66 18 68
rect 12 64 14 66
rect 16 64 18 66
rect 12 62 18 64
rect -85 58 -79 60
rect -118 54 -112 56
rect -118 52 -116 54
rect -114 52 -112 54
rect -173 47 -171 49
rect -169 47 -164 49
rect -262 33 -260 38
rect -252 36 -250 41
rect -242 36 -240 41
rect -222 32 -220 36
rect -173 45 -164 47
rect -148 47 -146 50
rect -166 42 -164 45
rect -156 42 -154 46
rect -148 45 -144 47
rect -146 42 -144 45
rect -139 42 -137 51
rect -118 50 -112 52
rect -108 54 -102 56
rect -108 52 -106 54
rect -104 52 -102 54
rect -108 50 -102 52
rect -118 45 -116 50
rect -105 45 -103 50
rect -98 45 -96 58
rect -81 57 -79 58
rect -70 57 -68 60
rect -54 57 -52 60
rect -81 55 -68 57
rect -62 55 -52 57
rect -44 56 -42 60
rect -34 57 -32 60
rect -78 47 -76 55
rect -62 51 -60 55
rect -69 49 -60 51
rect -48 54 -42 56
rect -48 52 -46 54
rect -44 52 -42 54
rect -48 50 -42 52
rect -38 55 -32 57
rect -38 53 -36 55
rect -34 53 -32 55
rect -38 51 -32 53
rect 28 58 30 70
rect 140 99 142 103
rect 228 99 230 103
rect 240 99 242 103
rect 252 99 254 103
rect 260 99 262 103
rect 272 99 274 103
rect 284 99 286 103
rect 292 99 294 103
rect 120 90 122 94
rect 128 90 130 94
rect 28 56 36 58
rect 28 54 32 56
rect 34 54 36 56
rect 28 52 36 54
rect -69 47 -67 49
rect -65 47 -60 49
rect -182 35 -180 38
rect -209 29 -207 34
rect -202 29 -200 34
rect -182 33 -177 35
rect -179 25 -177 33
rect -166 29 -164 33
rect -156 25 -154 33
rect -118 32 -116 36
rect -69 45 -60 47
rect -44 47 -42 50
rect -62 42 -60 45
rect -52 42 -50 46
rect -44 45 -40 47
rect -42 42 -40 45
rect -35 42 -33 51
rect 12 46 18 48
rect 12 44 14 46
rect 16 44 18 46
rect 12 42 18 44
rect 22 46 28 48
rect 40 46 42 60
rect 120 58 122 61
rect 116 56 122 58
rect 128 58 130 61
rect 216 75 218 79
rect 128 56 136 58
rect 116 48 118 56
rect 128 54 132 56
rect 134 54 136 56
rect 128 52 136 54
rect 22 44 24 46
rect 26 44 42 46
rect 22 42 28 44
rect -78 35 -76 38
rect -146 25 -144 30
rect -139 25 -137 30
rect -179 23 -154 25
rect -105 29 -103 34
rect -98 29 -96 34
rect -78 33 -73 35
rect -75 25 -73 33
rect -62 29 -60 33
rect -52 25 -50 33
rect 16 39 18 42
rect -42 25 -40 30
rect -35 25 -33 30
rect -75 23 -50 25
rect 28 36 36 38
rect 28 34 32 36
rect 34 34 36 36
rect 28 32 36 34
rect 28 29 30 32
rect 40 30 42 44
rect 112 46 118 48
rect 112 44 114 46
rect 116 44 118 46
rect 112 42 118 44
rect 122 46 128 48
rect 140 46 142 60
rect 216 58 218 61
rect 208 56 218 58
rect 208 54 210 56
rect 212 54 218 56
rect 208 52 218 54
rect 122 44 124 46
rect 126 44 142 46
rect 122 42 128 44
rect 116 30 118 42
rect 128 36 136 38
rect 128 34 132 36
rect 134 34 136 36
rect 128 32 136 34
rect 16 15 18 19
rect 128 29 130 32
rect 140 30 142 44
rect 216 42 218 52
rect 228 58 230 80
rect 240 78 242 81
rect 234 76 242 78
rect 234 74 236 76
rect 238 74 242 76
rect 234 72 242 74
rect 228 56 234 58
rect 228 54 230 56
rect 232 54 234 56
rect 228 52 234 54
rect 116 16 118 20
rect 128 15 130 19
rect 216 30 218 34
rect 228 28 230 52
rect 240 46 242 72
rect 252 68 254 80
rect 248 66 254 68
rect 248 64 250 66
rect 252 64 254 66
rect 248 62 254 64
rect 248 56 254 58
rect 260 56 262 80
rect 272 77 274 80
rect 284 77 286 80
rect 248 54 250 56
rect 252 54 262 56
rect 248 52 254 54
rect 240 44 254 46
rect 234 36 242 38
rect 234 34 236 36
rect 238 34 242 36
rect 234 32 242 34
rect 240 28 242 32
rect 252 28 254 44
rect 260 28 262 54
rect 270 75 274 77
rect 280 75 286 77
rect 270 38 272 75
rect 280 58 282 75
rect 292 68 294 80
rect 304 74 306 78
rect 286 66 294 68
rect 286 64 288 66
rect 290 64 294 66
rect 286 62 294 64
rect 276 56 282 58
rect 304 56 306 60
rect 276 54 278 56
rect 280 54 306 56
rect 276 52 282 54
rect 280 44 282 52
rect 266 36 272 38
rect 266 34 268 36
rect 270 34 272 36
rect 266 32 272 34
rect 276 42 282 44
rect 286 46 294 48
rect 286 44 288 46
rect 290 44 294 46
rect 286 42 294 44
rect 304 42 306 54
rect 276 28 278 42
rect 282 36 288 38
rect 282 34 284 36
rect 286 34 288 36
rect 282 32 288 34
rect 272 26 278 28
rect 272 23 274 26
rect 284 24 286 32
rect 292 24 294 42
rect 304 30 306 34
rect 228 12 230 16
rect 240 12 242 16
rect 252 12 254 16
rect 260 12 262 16
rect 28 7 30 11
rect 40 7 42 11
rect 140 7 142 11
rect 272 7 274 11
rect 284 8 286 12
rect 292 8 294 12
<< ndif >>
rect -269 45 -262 47
rect -269 43 -267 45
rect -265 43 -262 45
rect -269 41 -262 43
rect -267 38 -262 41
rect -260 41 -252 47
rect -250 45 -242 47
rect -250 43 -247 45
rect -245 43 -242 45
rect -250 41 -242 43
rect -240 41 -233 47
rect -189 45 -182 47
rect -227 42 -222 45
rect -260 38 -254 41
rect -258 34 -254 38
rect -238 34 -233 41
rect -229 40 -222 42
rect -229 38 -227 40
rect -225 38 -222 40
rect -229 36 -222 38
rect -220 36 -209 45
rect -258 32 -252 34
rect -258 30 -256 32
rect -254 30 -252 32
rect -258 28 -252 30
rect -239 32 -233 34
rect -218 34 -209 36
rect -207 34 -202 45
rect -200 40 -195 45
rect -189 43 -187 45
rect -185 43 -182 45
rect -189 41 -182 43
rect -200 38 -193 40
rect -187 38 -182 41
rect -180 42 -175 47
rect -85 45 -78 47
rect -123 42 -118 45
rect -180 38 -166 42
rect -200 36 -197 38
rect -195 36 -193 38
rect -200 34 -193 36
rect -175 37 -166 38
rect -175 35 -173 37
rect -171 35 -166 37
rect -239 30 -237 32
rect -235 30 -233 32
rect -239 28 -233 30
rect -218 28 -211 34
rect -175 33 -166 35
rect -164 40 -156 42
rect -164 38 -161 40
rect -159 38 -156 40
rect -164 33 -156 38
rect -154 38 -146 42
rect -154 36 -151 38
rect -149 36 -146 38
rect -154 33 -146 36
rect -218 26 -216 28
rect -214 26 -211 28
rect -218 24 -211 26
rect -151 30 -146 33
rect -144 30 -139 42
rect -137 30 -129 42
rect -125 40 -118 42
rect -125 38 -123 40
rect -121 38 -118 40
rect -125 36 -118 38
rect -116 36 -105 45
rect -114 34 -105 36
rect -103 34 -98 45
rect -96 40 -91 45
rect -85 43 -83 45
rect -81 43 -78 45
rect -85 41 -78 43
rect -96 38 -89 40
rect -83 38 -78 41
rect -76 42 -71 47
rect -76 38 -62 42
rect -96 36 -93 38
rect -91 36 -89 38
rect -96 34 -89 36
rect -71 37 -62 38
rect -71 35 -69 37
rect -67 35 -62 37
rect -135 28 -129 30
rect -135 26 -133 28
rect -131 26 -129 28
rect -135 24 -129 26
rect -114 28 -107 34
rect -71 33 -62 35
rect -60 40 -52 42
rect -60 38 -57 40
rect -55 38 -52 40
rect -60 33 -52 38
rect -50 38 -42 42
rect -50 36 -47 38
rect -45 36 -42 38
rect -50 33 -42 36
rect -114 26 -112 28
rect -110 26 -107 28
rect -114 24 -107 26
rect -47 30 -42 33
rect -40 30 -35 42
rect -33 30 -25 42
rect -31 28 -25 30
rect -31 26 -29 28
rect -27 26 -25 28
rect -31 24 -25 26
rect 8 26 16 39
rect 8 24 10 26
rect 12 24 16 26
rect 8 19 16 24
rect 18 29 26 39
rect 35 29 40 30
rect 18 19 28 29
rect 20 11 28 19
rect 30 16 40 29
rect 30 14 34 16
rect 36 14 40 16
rect 30 11 40 14
rect 42 26 50 30
rect 42 24 46 26
rect 48 24 50 26
rect 42 11 50 24
rect 108 20 116 30
rect 118 29 123 30
rect 208 34 216 42
rect 218 38 226 42
rect 218 36 222 38
rect 224 36 226 38
rect 218 34 226 36
rect 135 29 140 30
rect 118 26 128 29
rect 118 24 122 26
rect 124 24 128 26
rect 118 20 128 24
rect 108 16 114 20
rect 120 19 128 20
rect 130 19 140 29
rect 108 14 110 16
rect 112 14 114 16
rect 132 16 140 19
rect 108 12 114 14
rect 132 14 134 16
rect 136 14 140 16
rect 132 11 140 14
rect 142 26 150 30
rect 142 24 146 26
rect 148 24 150 26
rect 142 11 150 24
rect 208 26 214 34
rect 244 36 250 38
rect 244 34 246 36
rect 248 34 250 36
rect 244 28 250 34
rect 208 24 210 26
rect 212 24 214 26
rect 208 22 214 24
rect 220 26 228 28
rect 220 24 222 26
rect 224 24 228 26
rect 220 16 228 24
rect 230 16 240 28
rect 242 16 252 28
rect 254 16 260 28
rect 262 26 270 28
rect 262 24 266 26
rect 268 24 270 26
rect 262 23 270 24
rect 296 38 304 42
rect 296 36 298 38
rect 300 36 304 38
rect 296 34 304 36
rect 306 34 314 42
rect 296 26 302 28
rect 296 24 298 26
rect 300 24 302 26
rect 279 23 284 24
rect 262 16 272 23
rect 264 11 272 16
rect 274 16 284 23
rect 274 14 278 16
rect 280 14 284 16
rect 274 12 284 14
rect 286 12 292 24
rect 294 12 302 24
rect 308 16 314 34
rect 308 14 310 16
rect 312 14 314 16
rect 308 12 314 14
rect 274 11 281 12
<< pdif >>
rect 8 96 14 98
rect 8 94 10 96
rect 12 94 14 96
rect 32 96 40 99
rect 8 91 14 94
rect 32 94 34 96
rect 36 94 40 96
rect -258 85 -249 87
rect -258 83 -256 85
rect -254 83 -249 85
rect -258 77 -249 83
rect -269 75 -262 77
rect -269 73 -267 75
rect -265 73 -262 75
rect -269 68 -262 73
rect -269 66 -267 68
rect -265 66 -262 68
rect -269 59 -262 66
rect -260 66 -249 77
rect -247 66 -242 87
rect -240 80 -235 87
rect -240 78 -233 80
rect -218 78 -212 80
rect -240 76 -237 78
rect -235 76 -233 78
rect -240 74 -233 76
rect -240 66 -235 74
rect -227 73 -222 78
rect -229 71 -222 73
rect -229 69 -227 71
rect -225 69 -222 71
rect -260 59 -252 66
rect -229 64 -222 69
rect -229 62 -227 64
rect -225 62 -222 64
rect -229 60 -222 62
rect -220 76 -212 78
rect -220 74 -217 76
rect -215 74 -212 76
rect -220 67 -212 74
rect -210 78 -202 80
rect -210 76 -207 78
rect -205 76 -202 78
rect -210 71 -202 76
rect -210 69 -207 71
rect -205 69 -202 71
rect -210 67 -202 69
rect -200 78 -193 80
rect -200 76 -197 78
rect -195 76 -193 78
rect -200 67 -193 76
rect -220 60 -214 67
rect -179 66 -174 87
rect -181 64 -174 66
rect -181 62 -179 64
rect -177 62 -174 64
rect -181 60 -174 62
rect -172 85 -160 87
rect -172 83 -169 85
rect -167 83 -160 85
rect -172 78 -160 83
rect -143 78 -138 87
rect -172 76 -169 78
rect -167 76 -158 78
rect -172 60 -158 76
rect -156 71 -148 78
rect -156 69 -153 71
rect -151 69 -148 71
rect -156 64 -148 69
rect -156 62 -153 64
rect -151 62 -148 64
rect -156 60 -148 62
rect -146 71 -138 78
rect -146 69 -143 71
rect -141 69 -138 71
rect -146 60 -138 69
rect -136 81 -131 87
rect -136 79 -129 81
rect -136 77 -133 79
rect -131 77 -129 79
rect -114 78 -108 80
rect -136 75 -129 77
rect -136 60 -131 75
rect -123 73 -118 78
rect -125 71 -118 73
rect -125 69 -123 71
rect -121 69 -118 71
rect -125 64 -118 69
rect -125 62 -123 64
rect -121 62 -118 64
rect -125 60 -118 62
rect -116 76 -108 78
rect -116 74 -113 76
rect -111 74 -108 76
rect -116 67 -108 74
rect -106 78 -98 80
rect -106 76 -103 78
rect -101 76 -98 78
rect -106 71 -98 76
rect -106 69 -103 71
rect -101 69 -98 71
rect -106 67 -98 69
rect -96 78 -89 80
rect -96 76 -93 78
rect -91 76 -89 78
rect -96 67 -89 76
rect -116 60 -110 67
rect -75 66 -70 87
rect -77 64 -70 66
rect -77 62 -75 64
rect -73 62 -70 64
rect -77 60 -70 62
rect -68 85 -56 87
rect -68 83 -65 85
rect -63 83 -56 85
rect -68 78 -56 83
rect -39 78 -34 87
rect -68 76 -65 78
rect -63 76 -54 78
rect -68 60 -54 76
rect -52 71 -44 78
rect -52 69 -49 71
rect -47 69 -44 71
rect -52 64 -44 69
rect -52 62 -49 64
rect -47 62 -44 64
rect -52 60 -44 62
rect -42 71 -34 78
rect -42 69 -39 71
rect -37 69 -34 71
rect -42 60 -34 69
rect -32 81 -27 87
rect 8 86 16 91
rect 8 84 10 86
rect 12 84 16 86
rect -32 79 -25 81
rect -32 77 -29 79
rect -27 77 -25 79
rect -32 75 -25 77
rect -32 60 -27 75
rect 8 71 16 84
rect 18 90 26 91
rect 32 90 40 94
rect 18 86 28 90
rect 18 84 22 86
rect 24 84 28 86
rect 18 71 28 84
rect 23 70 28 71
rect 30 70 40 90
rect 32 60 40 70
rect 42 86 50 99
rect 132 96 140 99
rect 132 94 134 96
rect 136 94 140 96
rect 132 90 140 94
rect 42 84 46 86
rect 48 84 50 86
rect 42 76 50 84
rect 42 74 46 76
rect 48 74 50 76
rect 42 66 50 74
rect 42 64 46 66
rect 48 64 50 66
rect 42 60 50 64
rect 108 86 120 90
rect 108 84 110 86
rect 112 84 120 86
rect 108 61 120 84
rect 122 61 128 90
rect 130 61 140 90
rect 108 60 114 61
rect 135 60 140 61
rect 142 86 150 99
rect 142 84 146 86
rect 148 84 150 86
rect 142 76 150 84
rect 142 74 146 76
rect 148 74 150 76
rect 142 66 150 74
rect 142 64 146 66
rect 148 64 150 66
rect 142 60 150 64
rect 208 86 214 88
rect 208 84 210 86
rect 212 84 214 86
rect 208 75 214 84
rect 220 86 228 99
rect 220 84 222 86
rect 224 84 228 86
rect 220 80 228 84
rect 230 81 240 99
rect 242 81 252 99
rect 230 80 235 81
rect 208 61 216 75
rect 218 66 226 75
rect 218 64 222 66
rect 224 64 226 66
rect 218 61 226 64
rect 244 80 252 81
rect 254 80 260 99
rect 262 86 272 99
rect 262 84 266 86
rect 268 84 272 86
rect 262 80 272 84
rect 274 96 284 99
rect 274 94 278 96
rect 280 94 284 96
rect 274 80 284 94
rect 286 80 292 99
rect 294 86 302 99
rect 294 84 298 86
rect 300 84 302 86
rect 294 80 302 84
rect 308 86 314 88
rect 308 84 310 86
rect 312 84 314 86
rect 244 76 250 80
rect 244 74 246 76
rect 248 74 250 76
rect 244 72 250 74
rect 308 74 314 84
rect 296 66 304 74
rect 296 64 298 66
rect 300 64 304 66
rect 296 60 304 64
rect 306 60 314 74
<< alu1 >>
rect -273 100 323 105
rect -273 98 110 100
rect 112 98 122 100
rect 124 98 323 100
rect -273 96 323 98
rect -273 94 10 96
rect 12 94 34 96
rect 36 94 134 96
rect 136 94 278 96
rect 280 94 323 96
rect -273 93 323 94
rect -273 88 -21 93
rect -273 86 -266 88
rect -264 86 -226 88
rect -224 86 -153 88
rect -151 86 -122 88
rect -120 86 -49 88
rect -47 86 -21 88
rect -273 85 -21 86
rect 9 86 13 93
rect -269 79 -265 80
rect -269 75 -256 79
rect -269 73 -267 75
rect -269 68 -265 73
rect -269 66 -267 68
rect -269 56 -265 66
rect -237 67 -233 72
rect -269 54 -268 56
rect -266 54 -265 56
rect -269 47 -265 54
rect -237 65 -236 67
rect -234 65 -233 67
rect -237 63 -233 65
rect -254 61 -233 63
rect -254 59 -240 61
rect -238 59 -233 61
rect -229 71 -224 73
rect -229 69 -227 71
rect -225 69 -224 71
rect -189 74 -177 80
rect -229 67 -224 69
rect -229 65 -228 67
rect -226 65 -224 67
rect -229 64 -224 65
rect -229 62 -227 64
rect -225 62 -224 64
rect -229 60 -224 62
rect -197 69 -193 72
rect -197 67 -196 69
rect -194 67 -193 69
rect -269 45 -264 47
rect -269 43 -267 45
rect -265 43 -264 45
rect -269 41 -264 43
rect -254 54 -233 55
rect -254 52 -250 54
rect -248 52 -236 54
rect -234 52 -233 54
rect -254 51 -233 52
rect -237 42 -233 51
rect -229 40 -225 60
rect -197 63 -193 67
rect -206 62 -193 63
rect -206 60 -200 62
rect -198 60 -193 62
rect -206 59 -193 60
rect -189 69 -184 74
rect -189 67 -187 69
rect -185 67 -184 69
rect -189 62 -184 67
rect -189 60 -187 62
rect -185 60 -184 62
rect -189 58 -184 60
rect -214 54 -200 55
rect -214 52 -210 54
rect -208 52 -200 54
rect -214 51 -200 52
rect -229 38 -227 40
rect -225 38 -217 40
rect -229 34 -217 38
rect -205 45 -200 51
rect -205 43 -204 45
rect -202 43 -200 45
rect -205 42 -200 43
rect -173 49 -168 56
rect -145 71 -129 72
rect -145 69 -143 71
rect -141 69 -129 71
rect -145 67 -129 69
rect -133 62 -129 67
rect -133 60 -132 62
rect -130 60 -129 62
rect -173 48 -171 49
rect -181 47 -171 48
rect -169 47 -168 49
rect -181 45 -168 47
rect -181 43 -179 45
rect -177 43 -168 45
rect -181 42 -168 43
rect -133 39 -129 60
rect -153 38 -129 39
rect -153 36 -151 38
rect -149 36 -129 38
rect -153 35 -129 36
rect -125 71 -120 73
rect -125 69 -123 71
rect -121 69 -120 71
rect -85 74 -73 80
rect 9 84 10 86
rect 12 84 13 86
rect 9 82 13 84
rect 20 86 26 87
rect 20 84 22 86
rect 24 84 26 86
rect 20 83 26 84
rect -125 64 -120 69
rect -125 62 -123 64
rect -121 62 -120 64
rect -125 60 -120 62
rect -93 69 -89 72
rect -93 67 -92 69
rect -90 67 -89 69
rect -125 54 -121 60
rect -125 52 -124 54
rect -122 52 -121 54
rect -125 40 -121 52
rect -93 63 -89 67
rect -102 62 -89 63
rect -102 60 -101 62
rect -99 60 -96 62
rect -94 60 -89 62
rect -102 59 -89 60
rect -85 69 -80 74
rect -85 67 -83 69
rect -81 67 -80 69
rect -85 62 -80 67
rect -85 60 -83 62
rect -81 60 -80 62
rect -85 58 -80 60
rect -110 54 -96 55
rect -110 52 -106 54
rect -104 52 -96 54
rect -110 51 -96 52
rect -125 38 -123 40
rect -121 38 -113 40
rect -125 34 -113 38
rect -101 45 -96 51
rect -101 43 -100 45
rect -98 43 -96 45
rect -101 42 -96 43
rect -69 49 -64 56
rect -41 71 -25 72
rect -41 69 -39 71
rect -37 69 -25 71
rect -41 67 -25 69
rect -29 51 -25 67
rect 13 66 17 78
rect 13 64 14 66
rect 16 64 17 66
rect -69 48 -67 49
rect -77 47 -67 48
rect -65 47 -64 49
rect -77 45 -64 47
rect -77 43 -75 45
rect -73 43 -64 45
rect -77 42 -64 43
rect -29 50 -21 51
rect -29 48 -24 50
rect -22 48 -21 50
rect -29 47 -21 48
rect -29 39 -25 47
rect -49 38 -25 39
rect -49 36 -47 38
rect -45 36 -25 38
rect -49 35 -25 36
rect 13 46 17 64
rect 13 44 14 46
rect 16 44 17 46
rect 13 32 17 44
rect 22 47 26 83
rect 33 57 37 88
rect 30 56 37 57
rect 30 54 32 56
rect 34 54 37 56
rect 30 53 37 54
rect 22 46 28 47
rect 22 44 24 46
rect 26 44 28 46
rect 22 43 28 44
rect -273 28 -21 29
rect -273 26 -266 28
rect -264 26 -226 28
rect -224 26 -216 28
rect -214 26 -186 28
rect -184 26 -133 28
rect -131 26 -122 28
rect -120 26 -112 28
rect -110 26 -82 28
rect -80 26 -29 28
rect -27 26 -21 28
rect 22 27 26 43
rect 33 37 37 53
rect 30 36 37 37
rect 30 34 32 36
rect 34 34 37 36
rect 30 33 37 34
rect -273 17 -21 26
rect 8 26 26 27
rect 8 24 10 26
rect 12 24 26 26
rect 8 23 26 24
rect 33 22 37 33
rect 43 87 47 88
rect 43 86 50 87
rect 43 84 46 86
rect 48 84 50 86
rect 43 83 50 84
rect 108 86 126 87
rect 108 84 110 86
rect 112 84 126 86
rect 108 83 126 84
rect 43 77 47 83
rect 43 76 50 77
rect 43 74 46 76
rect 48 74 50 76
rect 43 73 50 74
rect 43 67 47 73
rect 43 66 50 67
rect 43 64 46 66
rect 48 64 50 66
rect 43 63 50 64
rect 43 57 47 63
rect 43 56 51 57
rect 43 54 48 56
rect 50 54 51 56
rect 43 53 51 54
rect 43 27 47 53
rect 113 46 117 78
rect 113 44 114 46
rect 116 44 117 46
rect 113 32 117 44
rect 122 47 126 83
rect 133 57 137 88
rect 130 56 137 57
rect 130 54 132 56
rect 134 54 137 56
rect 130 53 137 54
rect 122 46 128 47
rect 122 44 124 46
rect 126 44 128 46
rect 122 43 128 44
rect 122 27 126 43
rect 133 37 137 53
rect 130 36 137 37
rect 130 34 132 36
rect 134 34 137 36
rect 130 33 137 34
rect 43 26 50 27
rect 43 24 46 26
rect 48 24 50 26
rect 43 23 50 24
rect 120 26 126 27
rect 120 24 122 26
rect 124 24 126 26
rect 120 23 126 24
rect 43 22 47 23
rect 133 22 137 33
rect 143 87 147 88
rect 143 86 150 87
rect 143 84 146 86
rect 148 84 150 86
rect 143 83 150 84
rect 209 86 213 93
rect 209 84 210 86
rect 212 84 213 86
rect 143 77 147 83
rect 209 82 213 84
rect 220 86 270 87
rect 220 84 222 86
rect 224 84 266 86
rect 268 84 270 86
rect 220 83 270 84
rect 297 86 301 88
rect 297 84 298 86
rect 300 84 301 86
rect 209 77 213 78
rect 297 77 301 84
rect 309 86 313 93
rect 309 84 310 86
rect 312 84 313 86
rect 309 82 313 84
rect 309 77 313 78
rect 143 76 150 77
rect 143 74 146 76
rect 148 74 150 76
rect 143 73 150 74
rect 209 76 240 77
rect 209 74 236 76
rect 238 74 240 76
rect 209 73 240 74
rect 244 76 313 77
rect 244 74 246 76
rect 248 74 313 76
rect 244 73 313 74
rect 143 67 147 73
rect 143 66 150 67
rect 143 64 146 66
rect 148 64 150 66
rect 143 63 150 64
rect 143 57 147 63
rect 143 56 151 57
rect 143 54 148 56
rect 150 54 151 56
rect 143 53 151 54
rect 209 56 213 73
rect 209 54 210 56
rect 212 54 213 56
rect 143 27 147 53
rect 209 32 213 54
rect 219 66 254 67
rect 219 64 222 66
rect 224 64 250 66
rect 252 64 254 66
rect 219 63 254 64
rect 219 39 223 63
rect 229 56 233 58
rect 229 54 230 56
rect 232 54 233 56
rect 229 46 233 54
rect 240 56 254 57
rect 240 54 250 56
rect 252 54 254 56
rect 240 53 254 54
rect 259 47 263 73
rect 245 43 263 47
rect 269 57 273 68
rect 287 67 291 68
rect 278 66 291 67
rect 278 64 288 66
rect 290 64 291 66
rect 278 63 291 64
rect 296 66 303 67
rect 296 64 298 66
rect 300 64 303 66
rect 296 63 303 64
rect 287 57 291 63
rect 269 56 282 57
rect 269 54 278 56
rect 280 54 282 56
rect 269 53 282 54
rect 287 53 294 57
rect 219 38 226 39
rect 219 36 222 38
rect 224 37 226 38
rect 224 36 240 37
rect 219 34 236 36
rect 238 34 240 36
rect 219 33 240 34
rect 245 36 249 43
rect 269 42 273 53
rect 287 47 291 53
rect 278 46 291 47
rect 278 44 288 46
rect 290 44 291 46
rect 278 43 291 44
rect 287 42 291 43
rect 299 39 303 63
rect 296 38 303 39
rect 296 37 298 38
rect 245 34 246 36
rect 248 34 249 36
rect 245 32 249 34
rect 266 36 298 37
rect 300 36 303 38
rect 266 34 268 36
rect 270 34 284 36
rect 286 34 303 36
rect 266 33 303 34
rect 143 26 150 27
rect 143 24 146 26
rect 148 24 150 26
rect 143 23 150 24
rect 209 26 213 28
rect 309 27 313 73
rect 209 24 210 26
rect 212 24 213 26
rect 143 22 147 23
rect 209 17 213 24
rect 220 26 270 27
rect 220 24 222 26
rect 224 24 266 26
rect 268 24 270 26
rect 220 23 270 24
rect 296 26 313 27
rect 296 24 298 26
rect 300 24 313 26
rect 296 23 313 24
rect 309 22 313 23
rect -273 16 323 17
rect -273 14 34 16
rect 36 14 110 16
rect 112 14 134 16
rect 136 14 278 16
rect 280 14 310 16
rect 312 14 323 16
rect -273 5 323 14
<< alu2 >>
rect -275 95 196 99
rect -275 57 -271 95
rect -25 87 291 91
rect -197 69 -184 70
rect -237 67 -224 69
rect -237 65 -236 67
rect -234 65 -228 67
rect -226 65 -224 67
rect -197 67 -196 69
rect -194 67 -187 69
rect -185 67 -184 69
rect -197 66 -184 67
rect -93 69 -80 70
rect -93 67 -92 69
rect -90 67 -83 69
rect -81 67 -80 69
rect -93 66 -80 67
rect -237 64 -224 65
rect -133 62 -98 63
rect -133 60 -132 62
rect -130 60 -101 62
rect -99 60 -98 62
rect -133 59 -98 60
rect -275 56 -265 57
rect -275 54 -268 56
rect -266 54 -265 56
rect -275 53 -265 54
rect -237 54 -121 55
rect -237 52 -236 54
rect -234 52 -124 54
rect -122 52 -121 54
rect -237 51 -121 52
rect -25 51 -21 87
rect 51 79 253 83
rect 51 57 55 79
rect 155 71 233 75
rect 155 57 159 71
rect 47 56 55 57
rect 47 54 48 56
rect 50 54 55 56
rect 47 53 55 54
rect 147 56 159 57
rect 147 54 148 56
rect 150 54 159 56
rect 147 53 159 54
rect 229 56 233 71
rect 229 54 230 56
rect 232 54 233 56
rect 229 53 233 54
rect 249 56 253 79
rect 249 54 250 56
rect 252 54 253 56
rect 249 53 253 54
rect 287 66 291 87
rect 287 64 288 66
rect 290 64 291 66
rect -29 50 -21 51
rect -29 48 -24 50
rect -22 48 -21 50
rect -29 47 -21 48
rect -205 45 -173 47
rect -205 43 -204 45
rect -202 43 -179 45
rect -177 43 -173 45
rect -205 42 -173 43
rect -101 45 -69 47
rect -101 43 -100 45
rect -98 43 -75 45
rect -73 43 -69 45
rect 287 46 291 64
rect 287 44 288 46
rect 290 44 291 46
rect 287 43 291 44
rect -101 42 -69 43
<< ptie >>
rect -268 28 -262 30
rect -228 28 -222 30
rect -268 26 -266 28
rect -264 26 -262 28
rect -268 24 -262 26
rect -228 26 -226 28
rect -224 26 -222 28
rect -228 24 -222 26
rect -188 28 -182 30
rect -188 26 -186 28
rect -184 26 -182 28
rect -188 24 -182 26
rect -124 28 -118 30
rect -124 26 -122 28
rect -120 26 -118 28
rect -124 24 -118 26
rect -84 28 -78 30
rect -84 26 -82 28
rect -80 26 -78 28
rect -84 24 -78 26
<< ntie >>
rect 108 100 126 102
rect -268 88 -262 90
rect -268 86 -266 88
rect -264 86 -262 88
rect -228 88 -222 90
rect -268 84 -262 86
rect -228 86 -226 88
rect -224 86 -222 88
rect -155 88 -149 90
rect -228 84 -222 86
rect -155 86 -153 88
rect -151 86 -149 88
rect -124 88 -118 90
rect -155 84 -149 86
rect -124 86 -122 88
rect -120 86 -118 88
rect -51 88 -45 90
rect -124 84 -118 86
rect -51 86 -49 88
rect -47 86 -45 88
rect -51 84 -45 86
rect 108 98 110 100
rect 112 98 122 100
rect 124 98 126 100
rect 108 96 126 98
<< nmos >>
rect -262 38 -260 47
rect -252 41 -250 47
rect -242 41 -240 47
rect -222 36 -220 45
rect -209 34 -207 45
rect -202 34 -200 45
rect -182 38 -180 47
rect -166 33 -164 42
rect -156 33 -154 42
rect -146 30 -144 42
rect -139 30 -137 42
rect -118 36 -116 45
rect -105 34 -103 45
rect -98 34 -96 45
rect -78 38 -76 47
rect -62 33 -60 42
rect -52 33 -50 42
rect -42 30 -40 42
rect -35 30 -33 42
rect 16 19 18 39
rect 28 11 30 29
rect 40 11 42 30
rect 116 20 118 30
rect 216 34 218 42
rect 128 19 130 29
rect 140 11 142 30
rect 228 16 230 28
rect 240 16 242 28
rect 252 16 254 28
rect 260 16 262 28
rect 304 34 306 42
rect 272 11 274 23
rect 284 12 286 24
rect 292 12 294 24
<< pmos >>
rect -262 59 -260 77
rect -249 66 -247 87
rect -242 66 -240 87
rect -222 60 -220 78
rect -212 67 -210 80
rect -202 67 -200 80
rect -174 60 -172 87
rect -158 60 -156 78
rect -148 60 -146 78
rect -138 60 -136 87
rect -118 60 -116 78
rect -108 67 -106 80
rect -98 67 -96 80
rect -70 60 -68 87
rect -54 60 -52 78
rect -44 60 -42 78
rect -34 60 -32 87
rect 16 71 18 91
rect 28 70 30 90
rect 40 60 42 99
rect 120 61 122 90
rect 128 61 130 90
rect 140 60 142 99
rect 228 80 230 99
rect 240 81 242 99
rect 216 61 218 75
rect 252 80 254 99
rect 260 80 262 99
rect 272 80 274 99
rect 284 80 286 99
rect 292 80 294 99
rect 304 60 306 74
<< polyct0 >>
rect -260 52 -258 54
rect -220 52 -218 54
rect -150 52 -148 54
rect -140 53 -138 55
rect -116 52 -114 54
rect -46 52 -44 54
rect -36 53 -34 55
<< polyct1 >>
rect -240 59 -238 61
rect -250 52 -248 54
rect -200 60 -198 62
rect -187 60 -185 62
rect -210 52 -208 54
rect -96 60 -94 62
rect -83 60 -81 62
rect 14 64 16 66
rect -171 47 -169 49
rect -106 52 -104 54
rect 32 54 34 56
rect -67 47 -65 49
rect 14 44 16 46
rect 132 54 134 56
rect 24 44 26 46
rect 32 34 34 36
rect 114 44 116 46
rect 210 54 212 56
rect 124 44 126 46
rect 132 34 134 36
rect 236 74 238 76
rect 230 54 232 56
rect 250 64 252 66
rect 250 54 252 56
rect 236 34 238 36
rect 288 64 290 66
rect 278 54 280 56
rect 268 34 270 36
rect 288 44 290 46
rect 284 34 286 36
<< ndifct0 >>
rect -247 43 -245 45
rect -256 30 -254 32
rect -187 43 -185 45
rect -197 36 -195 38
rect -173 35 -171 37
rect -237 30 -235 32
rect -161 38 -159 40
rect -83 43 -81 45
rect -93 36 -91 38
rect -69 35 -67 37
rect -57 38 -55 40
<< ndifct1 >>
rect -267 43 -265 45
rect -227 38 -225 40
rect -151 36 -149 38
rect -216 26 -214 28
rect -123 38 -121 40
rect -133 26 -131 28
rect -47 36 -45 38
rect -112 26 -110 28
rect -29 26 -27 28
rect 10 24 12 26
rect 34 14 36 16
rect 46 24 48 26
rect 222 36 224 38
rect 122 24 124 26
rect 110 14 112 16
rect 134 14 136 16
rect 146 24 148 26
rect 246 34 248 36
rect 210 24 212 26
rect 222 24 224 26
rect 266 24 268 26
rect 298 36 300 38
rect 298 24 300 26
rect 278 14 280 16
rect 310 14 312 16
<< ntiect1 >>
rect -266 86 -264 88
rect -226 86 -224 88
rect -153 86 -151 88
rect -122 86 -120 88
rect -49 86 -47 88
rect 110 98 112 100
rect 122 98 124 100
<< ptiect1 >>
rect -266 26 -264 28
rect -226 26 -224 28
rect -186 26 -184 28
rect -122 26 -120 28
rect -82 26 -80 28
<< pdifct0 >>
rect -256 83 -254 85
rect -237 76 -235 78
rect -217 74 -215 76
rect -207 76 -205 78
rect -207 69 -205 71
rect -197 76 -195 78
rect -179 62 -177 64
rect -169 83 -167 85
rect -169 76 -167 78
rect -153 69 -151 71
rect -153 62 -151 64
rect -133 77 -131 79
rect -113 74 -111 76
rect -103 76 -101 78
rect -103 69 -101 71
rect -93 76 -91 78
rect -75 62 -73 64
rect -65 83 -63 85
rect -65 76 -63 78
rect -49 69 -47 71
rect -49 62 -47 64
rect -29 77 -27 79
<< pdifct1 >>
rect 10 94 12 96
rect 34 94 36 96
rect -267 73 -265 75
rect -267 66 -265 68
rect -227 69 -225 71
rect -227 62 -225 64
rect -143 69 -141 71
rect -123 69 -121 71
rect -123 62 -121 64
rect -39 69 -37 71
rect 10 84 12 86
rect 22 84 24 86
rect 134 94 136 96
rect 46 84 48 86
rect 46 74 48 76
rect 46 64 48 66
rect 110 84 112 86
rect 146 84 148 86
rect 146 74 148 76
rect 146 64 148 66
rect 210 84 212 86
rect 222 84 224 86
rect 222 64 224 66
rect 266 84 268 86
rect 278 94 280 96
rect 298 84 300 86
rect 310 84 312 86
rect 246 74 248 76
rect 298 64 300 66
<< alu0 >>
rect -258 83 -256 85
rect -254 83 -252 85
rect -258 82 -252 83
rect -250 78 -233 79
rect -250 76 -237 78
rect -235 76 -233 78
rect -250 75 -233 76
rect -219 76 -213 85
rect -265 64 -264 75
rect -250 71 -246 75
rect -219 74 -217 76
rect -215 74 -213 76
rect -219 73 -213 74
rect -208 78 -204 80
rect -208 76 -207 78
rect -205 76 -204 78
rect -261 67 -246 71
rect -261 54 -257 67
rect -208 71 -204 76
rect -199 78 -193 85
rect -170 83 -169 85
rect -167 83 -166 85
rect -199 76 -197 78
rect -195 76 -193 78
rect -199 75 -193 76
rect -170 78 -166 83
rect -170 76 -169 78
rect -167 76 -166 78
rect -170 74 -166 76
rect -162 79 -129 80
rect -162 77 -133 79
rect -131 77 -129 79
rect -162 76 -129 77
rect -115 76 -109 85
rect -208 70 -207 71
rect -221 69 -207 70
rect -205 69 -204 71
rect -221 66 -204 69
rect -242 58 -236 59
rect -261 52 -260 54
rect -258 52 -257 54
rect -261 46 -257 52
rect -261 45 -243 46
rect -261 43 -247 45
rect -245 43 -243 45
rect -261 42 -243 43
rect -221 54 -217 66
rect -162 65 -158 76
rect -115 74 -113 76
rect -111 74 -109 76
rect -115 73 -109 74
rect -104 78 -100 80
rect -104 76 -103 78
rect -101 76 -100 78
rect -181 64 -158 65
rect -181 62 -179 64
rect -177 62 -158 64
rect -181 61 -158 62
rect -181 55 -177 61
rect -221 52 -220 54
rect -218 52 -217 54
rect -221 47 -217 52
rect -221 43 -209 47
rect -225 40 -224 42
rect -213 39 -209 43
rect -188 51 -177 55
rect -188 45 -184 51
rect -162 55 -158 61
rect -154 71 -150 73
rect -154 69 -153 71
rect -151 69 -150 71
rect -154 64 -150 69
rect -154 62 -153 64
rect -151 63 -150 64
rect -151 62 -138 63
rect -154 59 -138 62
rect -142 57 -138 59
rect -142 55 -137 57
rect -162 54 -146 55
rect -162 52 -150 54
rect -148 52 -146 54
rect -162 51 -146 52
rect -142 53 -140 55
rect -138 53 -137 55
rect -142 51 -137 53
rect -188 43 -187 45
rect -185 43 -184 45
rect -188 41 -184 43
rect -142 47 -138 51
rect -162 43 -138 47
rect -162 40 -158 43
rect -213 38 -193 39
rect -162 38 -161 40
rect -159 38 -158 40
rect -213 36 -197 38
rect -195 36 -193 38
rect -213 35 -193 36
rect -175 37 -169 38
rect -175 35 -173 37
rect -171 35 -169 37
rect -162 36 -158 38
rect -104 71 -100 76
rect -95 78 -89 85
rect -66 83 -65 85
rect -63 83 -62 85
rect -95 76 -93 78
rect -91 76 -89 78
rect -95 75 -89 76
rect -66 78 -62 83
rect -66 76 -65 78
rect -63 76 -62 78
rect -66 74 -62 76
rect -58 79 -25 80
rect -58 77 -29 79
rect -27 77 -25 79
rect -58 76 -25 77
rect -104 70 -103 71
rect -117 69 -103 70
rect -101 69 -100 71
rect -117 66 -100 69
rect -117 54 -113 66
rect -58 65 -54 76
rect -77 64 -54 65
rect -77 62 -75 64
rect -73 62 -54 64
rect -77 61 -54 62
rect -77 55 -73 61
rect -117 52 -116 54
rect -114 52 -113 54
rect -117 47 -113 52
rect -117 43 -105 47
rect -121 40 -120 42
rect -258 32 -252 33
rect -258 30 -256 32
rect -254 30 -252 32
rect -258 29 -252 30
rect -239 32 -233 33
rect -239 30 -237 32
rect -235 30 -233 32
rect -239 29 -233 30
rect -175 29 -169 35
rect -109 39 -105 43
rect -84 51 -73 55
rect -84 45 -80 51
rect -58 55 -54 61
rect -50 71 -46 73
rect -50 69 -49 71
rect -47 69 -46 71
rect -50 64 -46 69
rect -50 62 -49 64
rect -47 63 -46 64
rect -47 62 -34 63
rect -50 59 -34 62
rect -38 57 -34 59
rect -38 55 -33 57
rect -58 54 -42 55
rect -58 52 -46 54
rect -44 52 -42 54
rect -58 51 -42 52
rect -38 53 -36 55
rect -34 53 -33 55
rect -38 51 -33 53
rect -84 43 -83 45
rect -81 43 -80 45
rect -84 41 -80 43
rect -38 47 -34 51
rect -58 43 -34 47
rect -58 40 -54 43
rect -109 38 -89 39
rect -58 38 -57 40
rect -55 38 -54 40
rect -109 36 -93 38
rect -91 36 -89 38
rect -109 35 -89 36
rect -71 37 -65 38
rect -71 35 -69 37
rect -67 35 -65 37
rect -58 36 -54 38
rect -71 29 -65 35
<< via1 >>
rect -268 54 -266 56
rect -236 65 -234 67
rect -228 65 -226 67
rect -196 67 -194 69
rect -236 52 -234 54
rect -187 67 -185 69
rect -204 43 -202 45
rect -132 60 -130 62
rect -179 43 -177 45
rect -92 67 -90 69
rect -124 52 -122 54
rect -101 60 -99 62
rect -83 67 -81 69
rect -100 43 -98 45
rect -75 43 -73 45
rect -24 48 -22 50
rect 48 54 50 56
rect 148 54 150 56
rect 230 54 232 56
rect 250 54 252 56
rect 288 64 290 66
rect 288 44 290 46
<< labels >>
rlabel alu1 30 11 30 11 6 vss
rlabel alu1 30 99 30 99 6 vdd
rlabel alu1 130 11 130 11 6 vss
rlabel alu1 130 99 130 99 6 vdd
rlabel alu1 15 55 15 55 1 a
rlabel alu1 35 55 35 55 1 b
rlabel alu1 45 55 45 55 1 andout
rlabel alu1 115 55 115 55 1 a
rlabel alu1 135 55 135 55 1 b
rlabel alu1 145 55 145 55 1 orout
rlabel polyct1 211 55 211 55 6 cmd1
rlabel polyct1 231 55 231 55 6 i2
rlabel alu1 221 75 221 75 6 cmd1
rlabel alu1 231 75 231 75 6 cmd1
rlabel alu1 261 11 261 11 6 vss
rlabel alu1 251 45 251 45 6 nq
rlabel polyct1 251 55 251 55 6 i1
rlabel alu1 261 55 261 55 6 nq
rlabel alu1 261 65 261 65 6 nq
rlabel alu1 251 75 251 75 6 nq
rlabel alu1 261 75 261 75 6 nq
rlabel alu1 261 99 261 99 6 vdd
rlabel alu1 281 45 281 45 6 i0
rlabel alu1 271 55 271 55 6 cmd0
rlabel alu1 291 55 291 55 6 i0
rlabel alu1 281 65 281 65 6 i0
rlabel alu1 271 75 271 75 6 nq
rlabel alu1 281 75 281 75 6 nq
rlabel alu1 291 75 291 75 6 nq
rlabel alu1 301 25 301 25 6 nq
rlabel alu1 311 50 311 50 6 nq
rlabel alu1 301 75 301 75 6 nq
rlabel alu0 -186 48 -186 48 6 bn
rlabel alu0 -140 53 -140 53 6 an
rlabel alu1 -171 49 -171 49 6 a
rlabel alu1 -159 25 -159 25 6 vss
rlabel alu1 -159 89 -159 89 6 vdd
rlabel alu1 -195 69 -195 69 6 b
rlabel alu1 -211 89 -211 89 6 vdd
rlabel alu1 -211 53 -211 53 6 a
rlabel alu1 -211 25 -211 25 6 vss
rlabel alu0 -219 56 -219 56 6 zn
rlabel alu1 -107 25 -107 25 6 vss
rlabel alu1 -107 89 -107 89 6 vdd
rlabel alu1 -27 49 -27 49 1 sum
rlabel alu1 -55 89 -55 89 6 vdd
rlabel alu1 -55 25 -55 25 6 vss
rlabel alu1 -131 49 -131 49 1 s
rlabel alu1 -107 52 -107 52 1 cin
rlabel alu1 -219 37 -219 37 1 co
rlabel alu0 -115 55 -115 55 1 zn_1
rlabel alu0 -82 48 -82 48 1 bn_1
rlabel alu0 -56 40 -56 40 1 an_1
rlabel alu1 -251 89 -251 89 6 vdd
rlabel alu1 -251 25 -251 25 6 vss
rlabel alu1 -115 37 -115 37 1 c1
rlabel alu0 -242 77 -242 77 1 zn_2
rlabel nwell -267 57 -267 57 1 cout
<< end >>
