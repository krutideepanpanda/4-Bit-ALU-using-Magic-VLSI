magic
tech scmos
timestamp 1636215170
<< ab >>
rect -25 91 223 93
rect -25 87 -8 91
rect -3 87 32 91
rect 36 87 85 91
rect 89 87 136 91
rect 140 87 189 91
rect 193 87 223 91
rect -25 85 223 87
rect -25 53 55 85
rect 56 53 159 85
rect 160 53 223 85
rect -25 27 223 53
rect -25 26 33 27
rect -25 23 -8 26
rect -4 23 33 26
rect 37 24 86 27
rect 88 26 189 27
rect 88 24 137 26
rect 37 23 137 24
rect -25 22 137 23
rect 141 24 189 26
rect 193 24 223 27
rect 141 22 223 24
rect -25 21 223 22
rect 232 91 272 93
rect 232 87 250 91
rect 254 87 272 91
rect 232 74 272 87
rect 232 72 246 74
rect 248 72 272 74
rect 232 57 272 72
rect 232 55 259 57
rect 261 55 272 57
rect 232 54 272 55
rect 232 52 267 54
rect 269 52 272 54
rect 232 38 272 52
rect 232 36 243 38
rect 245 36 259 38
rect 261 36 272 38
rect 232 27 272 36
rect 232 23 250 27
rect 254 23 272 27
rect 232 21 272 23
rect 280 91 320 93
rect 280 87 298 91
rect 302 87 320 91
rect 280 78 320 87
rect 280 76 290 78
rect 292 76 307 78
rect 309 76 320 78
rect 280 62 320 76
rect 280 60 315 62
rect 317 60 320 62
rect 280 57 320 60
rect 280 55 307 57
rect 309 55 320 57
rect 280 45 320 55
rect 280 43 300 45
rect 302 43 320 45
rect 280 26 320 43
rect 280 23 298 26
rect 302 23 320 26
rect 280 21 320 23
rect 329 90 393 93
rect 329 88 360 90
rect 362 88 393 90
rect 329 78 393 88
rect 329 76 340 78
rect 342 76 388 78
rect 390 76 393 78
rect 329 75 393 76
rect 329 72 355 75
rect 359 72 393 75
rect 329 70 393 72
rect 329 68 380 70
rect 382 68 393 70
rect 329 63 393 68
rect 329 62 376 63
rect 329 60 356 62
rect 358 61 376 62
rect 378 61 393 63
rect 358 60 393 61
rect 329 58 393 60
rect 329 56 340 58
rect 342 56 348 58
rect 350 56 393 58
rect 329 54 364 56
rect 366 54 393 56
rect 329 52 332 54
rect 334 52 372 54
rect 376 52 393 54
rect 329 51 393 52
rect 329 49 388 51
rect 390 49 393 51
rect 329 48 393 49
rect 329 46 360 48
rect 362 46 393 48
rect 329 44 380 46
rect 382 44 393 46
rect 329 38 393 44
rect 329 34 355 38
rect 357 34 393 38
rect 329 26 393 34
rect 329 24 360 26
rect 362 24 393 26
rect 329 21 393 24
rect 403 90 467 93
rect 403 88 434 90
rect 436 88 467 90
rect 403 78 467 88
rect 403 76 414 78
rect 416 76 462 78
rect 464 76 467 78
rect 403 75 467 76
rect 403 72 429 75
rect 433 72 467 75
rect 403 70 467 72
rect 403 68 454 70
rect 456 68 467 70
rect 403 63 467 68
rect 403 62 450 63
rect 403 60 430 62
rect 432 61 450 62
rect 452 61 467 63
rect 432 60 467 61
rect 403 58 467 60
rect 403 56 414 58
rect 416 56 422 58
rect 424 56 467 58
rect 403 54 438 56
rect 440 54 467 56
rect 403 52 406 54
rect 408 52 446 54
rect 448 52 467 54
rect 403 51 467 52
rect 403 49 462 51
rect 464 49 467 51
rect 403 48 467 49
rect 403 46 434 48
rect 436 46 467 48
rect 403 44 454 46
rect 456 44 467 46
rect 403 38 467 44
rect 403 34 429 38
rect 431 34 467 38
rect 403 26 467 34
rect 403 24 434 26
rect 436 24 467 26
rect 403 21 467 24
rect 477 90 541 93
rect 477 88 508 90
rect 510 88 541 90
rect 477 78 541 88
rect 477 76 488 78
rect 490 76 536 78
rect 538 76 541 78
rect 477 75 541 76
rect 477 72 503 75
rect 507 72 541 75
rect 477 70 541 72
rect 477 68 528 70
rect 530 68 541 70
rect 477 63 541 68
rect 477 62 524 63
rect 477 60 504 62
rect 506 61 524 62
rect 526 61 541 63
rect 506 60 541 61
rect 477 58 541 60
rect 477 57 488 58
rect 477 55 480 57
rect 482 56 488 57
rect 490 56 496 58
rect 498 56 541 58
rect 482 55 512 56
rect 477 54 512 55
rect 514 54 541 56
rect 477 52 480 54
rect 482 52 520 54
rect 522 52 541 54
rect 477 51 541 52
rect 477 49 536 51
rect 538 49 541 51
rect 477 48 541 49
rect 477 46 508 48
rect 510 46 541 48
rect 477 44 528 46
rect 530 44 541 46
rect 477 38 541 44
rect 477 34 503 38
rect 505 34 541 38
rect 477 26 541 34
rect 477 24 508 26
rect 510 24 541 26
rect 477 21 541 24
rect 50 16 56 21
rect 154 16 160 21
<< nwell >>
rect -30 53 546 98
<< pwell >>
rect -30 16 546 53
<< poly >>
rect -3 87 -1 91
rect 4 87 6 91
rect -16 77 -14 82
rect 72 87 74 91
rect 24 78 26 82
rect 34 80 36 85
rect 44 80 46 85
rect -16 56 -14 59
rect -3 56 -1 66
rect 4 63 6 66
rect 4 61 10 63
rect 4 59 6 61
rect 8 59 10 61
rect 4 57 10 59
rect -16 54 -10 56
rect -16 52 -14 54
rect -12 52 -10 54
rect -16 50 -10 52
rect -6 54 0 56
rect -6 52 -4 54
rect -2 52 0 54
rect -6 50 0 52
rect -16 47 -14 50
rect -6 47 -4 50
rect 4 47 6 57
rect 24 56 26 60
rect 34 56 36 67
rect 44 64 46 67
rect 44 62 50 64
rect 44 60 46 62
rect 48 60 50 62
rect 44 58 50 60
rect 57 62 63 64
rect 57 60 59 62
rect 61 60 63 62
rect 108 87 110 91
rect 88 78 90 82
rect 98 78 100 82
rect 176 87 178 91
rect 128 78 130 82
rect 138 80 140 85
rect 148 80 150 85
rect 57 58 63 60
rect 24 54 30 56
rect 24 52 26 54
rect 28 52 30 54
rect 24 50 30 52
rect 34 54 40 56
rect 34 52 36 54
rect 38 52 40 54
rect 34 50 40 52
rect 24 45 26 50
rect 37 45 39 50
rect 44 45 46 58
rect 61 57 63 58
rect 72 57 74 60
rect 88 57 90 60
rect 61 55 74 57
rect 80 55 90 57
rect 98 56 100 60
rect 108 57 110 60
rect 64 47 66 55
rect 80 51 82 55
rect 73 49 82 51
rect 94 54 100 56
rect 94 52 96 54
rect 98 52 100 54
rect 94 50 100 52
rect 104 55 110 57
rect 104 53 106 55
rect 108 53 110 55
rect 104 51 110 53
rect 128 56 130 60
rect 138 56 140 67
rect 148 64 150 67
rect 148 62 154 64
rect 148 60 150 62
rect 152 60 154 62
rect 148 58 154 60
rect 161 62 167 64
rect 161 60 163 62
rect 165 60 167 62
rect 212 87 214 91
rect 192 78 194 82
rect 202 78 204 82
rect 289 87 291 91
rect 296 87 298 91
rect 241 80 243 85
rect 251 80 253 85
rect 261 78 263 82
rect 241 64 243 67
rect 237 62 243 64
rect 237 60 239 62
rect 241 60 243 62
rect 161 58 167 60
rect 128 54 134 56
rect 128 52 130 54
rect 132 52 134 54
rect 73 47 75 49
rect 77 47 82 49
rect -16 33 -14 38
rect -6 36 -4 41
rect 4 36 6 41
rect 24 32 26 36
rect 73 45 82 47
rect 98 47 100 50
rect 80 42 82 45
rect 90 42 92 46
rect 98 45 102 47
rect 100 42 102 45
rect 107 42 109 51
rect 128 50 134 52
rect 138 54 144 56
rect 138 52 140 54
rect 142 52 144 54
rect 138 50 144 52
rect 128 45 130 50
rect 141 45 143 50
rect 148 45 150 58
rect 165 57 167 58
rect 176 57 178 60
rect 192 57 194 60
rect 165 55 178 57
rect 184 55 194 57
rect 202 56 204 60
rect 212 57 214 60
rect 237 58 243 60
rect 168 47 170 55
rect 184 51 186 55
rect 177 49 186 51
rect 198 54 204 56
rect 198 52 200 54
rect 202 52 204 54
rect 198 50 204 52
rect 208 55 214 57
rect 208 53 210 55
rect 212 53 214 55
rect 208 51 214 53
rect 177 47 179 49
rect 181 47 186 49
rect 64 35 66 38
rect 37 29 39 34
rect 44 29 46 34
rect 64 33 69 35
rect 67 25 69 33
rect 80 29 82 33
rect 90 25 92 33
rect 128 32 130 36
rect 177 45 186 47
rect 202 47 204 50
rect 184 42 186 45
rect 194 42 196 46
rect 202 45 206 47
rect 204 42 206 45
rect 211 42 213 51
rect 241 45 243 58
rect 251 56 253 67
rect 338 87 340 91
rect 348 87 350 91
rect 355 87 357 91
rect 365 87 367 91
rect 372 87 374 91
rect 412 87 414 91
rect 422 87 424 91
rect 429 87 431 91
rect 439 87 441 91
rect 446 87 448 91
rect 486 87 488 91
rect 496 87 498 91
rect 503 87 505 91
rect 513 87 515 91
rect 520 87 522 91
rect 309 77 311 82
rect 289 63 291 66
rect 285 61 291 63
rect 261 56 263 60
rect 285 59 287 61
rect 289 59 291 61
rect 285 57 291 59
rect 247 54 253 56
rect 247 52 249 54
rect 251 52 253 54
rect 247 50 253 52
rect 257 54 263 56
rect 257 52 259 54
rect 261 52 263 54
rect 257 50 263 52
rect 248 45 250 50
rect 261 45 263 50
rect 289 47 291 57
rect 296 56 298 66
rect 385 74 391 76
rect 385 72 387 74
rect 389 72 391 74
rect 309 56 311 59
rect 295 54 301 56
rect 295 52 297 54
rect 299 52 301 54
rect 295 50 301 52
rect 305 54 311 56
rect 305 52 307 54
rect 309 52 311 54
rect 305 50 311 52
rect 338 51 340 69
rect 348 61 350 71
rect 345 59 351 61
rect 345 57 347 59
rect 349 57 351 59
rect 345 55 351 57
rect 355 56 357 71
rect 365 66 367 71
rect 362 64 368 66
rect 362 62 364 64
rect 366 62 368 64
rect 362 60 368 62
rect 372 56 374 71
rect 382 70 391 72
rect 382 67 384 70
rect 459 74 465 76
rect 459 72 461 74
rect 463 72 465 74
rect 299 47 301 50
rect 309 47 311 50
rect 337 49 343 51
rect 337 47 339 49
rect 341 47 343 49
rect 168 35 170 38
rect 100 25 102 30
rect 107 25 109 30
rect 67 23 92 25
rect 141 29 143 34
rect 148 29 150 34
rect 168 33 173 35
rect 171 25 173 33
rect 184 29 186 33
rect 194 25 196 33
rect 204 25 206 30
rect 211 25 213 30
rect 241 29 243 34
rect 248 29 250 34
rect 171 23 196 25
rect 261 32 263 36
rect 289 36 291 41
rect 299 36 301 41
rect 337 45 343 47
rect 338 42 340 45
rect 309 33 311 38
rect 348 41 350 55
rect 355 54 367 56
rect 355 48 361 50
rect 355 46 357 48
rect 359 46 361 48
rect 355 44 361 46
rect 355 41 357 44
rect 365 41 367 54
rect 372 49 378 56
rect 372 47 374 49
rect 376 47 378 49
rect 372 45 378 47
rect 372 41 374 45
rect 382 41 384 59
rect 412 51 414 69
rect 422 61 424 71
rect 419 59 425 61
rect 419 57 421 59
rect 423 57 425 59
rect 419 55 425 57
rect 429 56 431 71
rect 439 66 441 71
rect 436 64 442 66
rect 436 62 438 64
rect 440 62 442 64
rect 436 60 442 62
rect 446 56 448 71
rect 456 70 465 72
rect 456 67 458 70
rect 533 74 539 76
rect 533 72 535 74
rect 537 72 539 74
rect 411 49 417 51
rect 411 47 413 49
rect 415 47 417 49
rect 411 45 417 47
rect 412 42 414 45
rect 338 28 340 33
rect 348 28 350 33
rect 355 28 357 33
rect 365 25 367 33
rect 372 29 374 33
rect 382 25 384 35
rect 422 41 424 55
rect 429 54 441 56
rect 429 48 435 50
rect 429 46 431 48
rect 433 46 435 48
rect 429 44 435 46
rect 429 41 431 44
rect 439 41 441 54
rect 446 54 452 56
rect 446 52 448 54
rect 450 52 452 54
rect 446 50 452 52
rect 446 41 448 50
rect 456 41 458 59
rect 486 51 488 69
rect 496 61 498 71
rect 493 59 499 61
rect 493 57 495 59
rect 497 57 499 59
rect 493 55 499 57
rect 503 56 505 71
rect 513 66 515 71
rect 510 64 516 66
rect 510 62 512 64
rect 514 62 516 64
rect 510 60 516 62
rect 520 56 522 71
rect 530 70 539 72
rect 530 67 532 70
rect 485 49 491 51
rect 485 47 487 49
rect 489 47 491 49
rect 485 45 491 47
rect 486 42 488 45
rect 412 28 414 33
rect 422 28 424 33
rect 429 28 431 33
rect 365 23 384 25
rect 439 25 441 33
rect 446 29 448 33
rect 456 25 458 35
rect 496 41 498 55
rect 503 54 515 56
rect 503 48 509 50
rect 503 46 505 48
rect 507 46 509 48
rect 503 44 509 46
rect 503 41 505 44
rect 513 41 515 54
rect 520 54 526 56
rect 520 52 522 54
rect 524 52 526 54
rect 520 50 526 52
rect 520 41 522 50
rect 530 41 532 59
rect 486 28 488 33
rect 496 28 498 33
rect 503 28 505 33
rect 439 23 458 25
rect 513 25 515 33
rect 520 29 522 33
rect 530 25 532 35
rect 513 23 532 25
<< ndif >>
rect -23 45 -16 47
rect -23 43 -21 45
rect -19 43 -16 45
rect -23 41 -16 43
rect -21 38 -16 41
rect -14 41 -6 47
rect -4 45 4 47
rect -4 43 -1 45
rect 1 43 4 45
rect -4 41 4 43
rect 6 41 13 47
rect 57 45 64 47
rect 19 42 24 45
rect -14 38 -8 41
rect -12 34 -8 38
rect 8 34 13 41
rect 17 40 24 42
rect 17 38 19 40
rect 21 38 24 40
rect 17 36 24 38
rect 26 36 37 45
rect -12 32 -6 34
rect -12 30 -10 32
rect -8 30 -6 32
rect -12 28 -6 30
rect 7 32 13 34
rect 28 34 37 36
rect 39 34 44 45
rect 46 40 51 45
rect 57 43 59 45
rect 61 43 64 45
rect 57 41 64 43
rect 46 38 53 40
rect 59 38 64 41
rect 66 42 71 47
rect 161 45 168 47
rect 123 42 128 45
rect 66 38 80 42
rect 46 36 49 38
rect 51 36 53 38
rect 46 34 53 36
rect 71 37 80 38
rect 71 35 73 37
rect 75 35 80 37
rect 7 30 9 32
rect 11 30 13 32
rect 7 28 13 30
rect 28 28 35 34
rect 71 33 80 35
rect 82 40 90 42
rect 82 38 85 40
rect 87 38 90 40
rect 82 33 90 38
rect 92 38 100 42
rect 92 36 95 38
rect 97 36 100 38
rect 92 33 100 36
rect 28 26 30 28
rect 32 26 35 28
rect 28 24 35 26
rect 95 30 100 33
rect 102 30 107 42
rect 109 30 117 42
rect 121 40 128 42
rect 121 38 123 40
rect 125 38 128 40
rect 121 36 128 38
rect 130 36 141 45
rect 132 34 141 36
rect 143 34 148 45
rect 150 40 155 45
rect 161 43 163 45
rect 165 43 168 45
rect 161 41 168 43
rect 150 38 157 40
rect 163 38 168 41
rect 170 42 175 47
rect 170 38 184 42
rect 150 36 153 38
rect 155 36 157 38
rect 150 34 157 36
rect 175 37 184 38
rect 175 35 177 37
rect 179 35 184 37
rect 111 28 117 30
rect 111 26 113 28
rect 115 26 117 28
rect 111 24 117 26
rect 132 28 139 34
rect 175 33 184 35
rect 186 40 194 42
rect 186 38 189 40
rect 191 38 194 40
rect 186 33 194 38
rect 196 38 204 42
rect 196 36 199 38
rect 201 36 204 38
rect 196 33 204 36
rect 132 26 134 28
rect 136 26 139 28
rect 132 24 139 26
rect 199 30 204 33
rect 206 30 211 42
rect 213 30 221 42
rect 236 40 241 45
rect 234 38 241 40
rect 234 36 236 38
rect 238 36 241 38
rect 234 34 241 36
rect 243 34 248 45
rect 250 36 261 45
rect 263 42 268 45
rect 263 40 270 42
rect 263 38 266 40
rect 268 38 270 40
rect 263 36 270 38
rect 282 41 289 47
rect 291 45 299 47
rect 291 43 294 45
rect 296 43 299 45
rect 291 41 299 43
rect 301 41 309 47
rect 250 34 259 36
rect 215 28 221 30
rect 215 26 217 28
rect 219 26 221 28
rect 215 24 221 26
rect 252 28 259 34
rect 282 34 287 41
rect 303 38 309 41
rect 311 45 318 47
rect 311 43 314 45
rect 316 43 318 45
rect 311 41 318 43
rect 311 38 316 41
rect 331 40 338 42
rect 331 38 333 40
rect 335 38 338 40
rect 303 34 307 38
rect 282 32 288 34
rect 282 30 284 32
rect 286 30 288 32
rect 252 26 255 28
rect 257 26 259 28
rect 252 24 259 26
rect 282 28 288 30
rect 301 32 307 34
rect 331 36 338 38
rect 333 33 338 36
rect 340 41 345 42
rect 340 37 348 41
rect 340 35 343 37
rect 345 35 348 37
rect 340 33 348 35
rect 350 33 355 41
rect 357 37 365 41
rect 357 35 360 37
rect 362 35 365 37
rect 357 33 365 35
rect 367 33 372 41
rect 374 39 382 41
rect 374 37 377 39
rect 379 37 382 39
rect 374 35 382 37
rect 384 39 391 41
rect 384 37 387 39
rect 389 37 391 39
rect 384 35 391 37
rect 405 40 412 42
rect 405 38 407 40
rect 409 38 412 40
rect 405 36 412 38
rect 374 33 380 35
rect 301 30 303 32
rect 305 30 307 32
rect 301 28 307 30
rect 407 33 412 36
rect 414 41 419 42
rect 414 37 422 41
rect 414 35 417 37
rect 419 35 422 37
rect 414 33 422 35
rect 424 33 429 41
rect 431 37 439 41
rect 431 35 434 37
rect 436 35 439 37
rect 431 33 439 35
rect 441 33 446 41
rect 448 39 456 41
rect 448 37 451 39
rect 453 37 456 39
rect 448 35 456 37
rect 458 39 465 41
rect 458 37 461 39
rect 463 37 465 39
rect 458 35 465 37
rect 479 40 486 42
rect 479 38 481 40
rect 483 38 486 40
rect 479 36 486 38
rect 448 33 454 35
rect 481 33 486 36
rect 488 41 493 42
rect 488 37 496 41
rect 488 35 491 37
rect 493 35 496 37
rect 488 33 496 35
rect 498 33 503 41
rect 505 37 513 41
rect 505 35 508 37
rect 510 35 513 37
rect 505 33 513 35
rect 515 33 520 41
rect 522 39 530 41
rect 522 37 525 39
rect 527 37 530 39
rect 522 35 530 37
rect 532 39 539 41
rect 532 37 535 39
rect 537 37 539 39
rect 532 35 539 37
rect 522 33 528 35
<< pdif >>
rect -12 85 -3 87
rect -12 83 -10 85
rect -8 83 -3 85
rect -12 77 -3 83
rect -23 75 -16 77
rect -23 73 -21 75
rect -19 73 -16 75
rect -23 68 -16 73
rect -23 66 -21 68
rect -19 66 -16 68
rect -23 64 -16 66
rect -21 59 -16 64
rect -14 66 -3 77
rect -1 66 4 87
rect 6 80 11 87
rect 6 78 13 80
rect 28 78 34 80
rect 6 76 9 78
rect 11 76 13 78
rect 6 74 13 76
rect 6 66 11 74
rect 19 73 24 78
rect 17 71 24 73
rect 17 69 19 71
rect 21 69 24 71
rect -14 59 -6 66
rect 17 64 24 69
rect 17 62 19 64
rect 21 62 24 64
rect 17 60 24 62
rect 26 76 34 78
rect 26 74 29 76
rect 31 74 34 76
rect 26 67 34 74
rect 36 78 44 80
rect 36 76 39 78
rect 41 76 44 78
rect 36 71 44 76
rect 36 69 39 71
rect 41 69 44 71
rect 36 67 44 69
rect 46 78 53 80
rect 46 76 49 78
rect 51 76 53 78
rect 46 67 53 76
rect 26 60 32 67
rect 67 66 72 87
rect 65 64 72 66
rect 65 62 67 64
rect 69 62 72 64
rect 65 60 72 62
rect 74 85 86 87
rect 74 83 77 85
rect 79 83 86 85
rect 74 78 86 83
rect 103 78 108 87
rect 74 76 77 78
rect 79 76 88 78
rect 74 60 88 76
rect 90 71 98 78
rect 90 69 93 71
rect 95 69 98 71
rect 90 64 98 69
rect 90 62 93 64
rect 95 62 98 64
rect 90 60 98 62
rect 100 71 108 78
rect 100 69 103 71
rect 105 69 108 71
rect 100 60 108 69
rect 110 81 115 87
rect 110 79 117 81
rect 110 77 113 79
rect 115 77 117 79
rect 132 78 138 80
rect 110 75 117 77
rect 110 60 115 75
rect 123 73 128 78
rect 121 71 128 73
rect 121 69 123 71
rect 125 69 128 71
rect 121 64 128 69
rect 121 62 123 64
rect 125 62 128 64
rect 121 60 128 62
rect 130 76 138 78
rect 130 74 133 76
rect 135 74 138 76
rect 130 67 138 74
rect 140 78 148 80
rect 140 76 143 78
rect 145 76 148 78
rect 140 71 148 76
rect 140 69 143 71
rect 145 69 148 71
rect 140 67 148 69
rect 150 78 157 80
rect 150 76 153 78
rect 155 76 157 78
rect 150 67 157 76
rect 130 60 136 67
rect 171 66 176 87
rect 169 64 176 66
rect 169 62 171 64
rect 173 62 176 64
rect 169 60 176 62
rect 178 85 190 87
rect 178 83 181 85
rect 183 83 190 85
rect 178 78 190 83
rect 207 78 212 87
rect 178 76 181 78
rect 183 76 192 78
rect 178 60 192 76
rect 194 71 202 78
rect 194 69 197 71
rect 199 69 202 71
rect 194 64 202 69
rect 194 62 197 64
rect 199 62 202 64
rect 194 60 202 62
rect 204 71 212 78
rect 204 69 207 71
rect 209 69 212 71
rect 204 60 212 69
rect 214 81 219 87
rect 214 79 221 81
rect 214 77 217 79
rect 219 77 221 79
rect 214 75 221 77
rect 234 78 241 80
rect 234 76 236 78
rect 238 76 241 78
rect 214 60 219 75
rect 234 67 241 76
rect 243 78 251 80
rect 243 76 246 78
rect 248 76 251 78
rect 243 71 251 76
rect 243 69 246 71
rect 248 69 251 71
rect 243 67 251 69
rect 253 78 259 80
rect 284 80 289 87
rect 282 78 289 80
rect 253 76 261 78
rect 253 74 256 76
rect 258 74 261 76
rect 253 67 261 74
rect 255 60 261 67
rect 263 73 268 78
rect 282 76 284 78
rect 286 76 289 78
rect 282 74 289 76
rect 263 71 270 73
rect 263 69 266 71
rect 268 69 270 71
rect 263 64 270 69
rect 284 66 289 74
rect 291 66 296 87
rect 298 85 307 87
rect 298 83 303 85
rect 305 83 307 85
rect 298 77 307 83
rect 333 80 338 87
rect 331 78 338 80
rect 298 66 309 77
rect 263 62 266 64
rect 268 62 270 64
rect 263 60 270 62
rect 301 59 309 66
rect 311 75 318 77
rect 311 73 314 75
rect 316 73 318 75
rect 331 76 333 78
rect 335 76 338 78
rect 331 74 338 76
rect 311 68 318 73
rect 333 69 338 74
rect 340 85 348 87
rect 340 83 343 85
rect 345 83 348 85
rect 340 71 348 83
rect 350 71 355 87
rect 357 75 365 87
rect 357 73 360 75
rect 362 73 365 75
rect 357 71 365 73
rect 367 71 372 87
rect 374 85 381 87
rect 374 83 377 85
rect 379 83 381 85
rect 374 75 381 83
rect 407 80 412 87
rect 405 78 412 80
rect 405 76 407 78
rect 409 76 412 78
rect 374 71 380 75
rect 405 74 412 76
rect 340 69 345 71
rect 311 66 314 68
rect 316 66 318 68
rect 311 64 318 66
rect 311 59 316 64
rect 376 67 380 71
rect 407 69 412 74
rect 414 85 422 87
rect 414 83 417 85
rect 419 83 422 85
rect 414 71 422 83
rect 424 71 429 87
rect 431 75 439 87
rect 431 73 434 75
rect 436 73 439 75
rect 431 71 439 73
rect 441 71 446 87
rect 448 85 455 87
rect 448 83 451 85
rect 453 83 455 85
rect 448 75 455 83
rect 481 80 486 87
rect 479 78 486 80
rect 479 76 481 78
rect 483 76 486 78
rect 448 71 454 75
rect 479 74 486 76
rect 414 69 419 71
rect 376 59 382 67
rect 384 65 389 67
rect 384 63 391 65
rect 384 61 387 63
rect 389 61 391 63
rect 384 59 391 61
rect 450 67 454 71
rect 481 69 486 74
rect 488 85 496 87
rect 488 83 491 85
rect 493 83 496 85
rect 488 71 496 83
rect 498 71 503 87
rect 505 75 513 87
rect 505 73 508 75
rect 510 73 513 75
rect 505 71 513 73
rect 515 71 520 87
rect 522 85 529 87
rect 522 83 525 85
rect 527 83 529 85
rect 522 75 529 83
rect 522 71 528 75
rect 488 69 493 71
rect 450 59 456 67
rect 458 65 463 67
rect 458 63 465 65
rect 458 61 461 63
rect 463 61 465 63
rect 458 59 465 61
rect 524 67 528 71
rect 524 59 530 67
rect 532 65 537 67
rect 532 63 539 65
rect 532 61 535 63
rect 537 61 539 63
rect 532 59 539 61
<< alu1 >>
rect -27 88 543 93
rect -27 86 -20 88
rect -18 86 20 88
rect 22 86 93 88
rect 95 86 124 88
rect 126 86 197 88
rect 199 86 265 88
rect 267 86 313 88
rect 315 86 543 88
rect -27 85 543 86
rect -23 79 -19 80
rect -23 75 -10 79
rect -23 73 -21 75
rect -23 68 -19 73
rect -23 66 -21 68
rect -23 47 -19 66
rect 9 67 13 72
rect 9 65 10 67
rect 12 65 13 67
rect 9 63 13 65
rect -8 61 13 63
rect -8 59 6 61
rect 8 59 13 61
rect 17 71 22 73
rect 17 69 19 71
rect 21 69 22 71
rect 57 74 69 80
rect 17 67 22 69
rect 17 65 18 67
rect 20 65 22 67
rect 17 64 22 65
rect 17 62 19 64
rect 21 62 22 64
rect 17 60 22 62
rect 49 69 53 72
rect 49 67 50 69
rect 52 67 53 69
rect -23 45 -18 47
rect -23 43 -21 45
rect -19 43 -18 45
rect -23 41 -18 43
rect -8 54 13 55
rect -8 52 -4 54
rect -2 52 10 54
rect 12 52 13 54
rect -8 51 13 52
rect 9 42 13 51
rect 17 40 21 60
rect 49 63 53 67
rect 40 62 53 63
rect 40 60 46 62
rect 48 60 53 62
rect 40 59 53 60
rect 57 69 62 74
rect 57 67 59 69
rect 61 67 62 69
rect 57 62 62 67
rect 57 60 59 62
rect 61 60 62 62
rect 57 58 62 60
rect 32 54 46 55
rect 32 52 36 54
rect 38 52 46 54
rect 32 51 46 52
rect 17 38 19 40
rect 21 38 29 40
rect 17 34 29 38
rect 41 45 46 51
rect 41 43 42 45
rect 44 43 46 45
rect 41 42 46 43
rect 73 49 78 56
rect 101 71 117 72
rect 101 69 103 71
rect 105 69 117 71
rect 101 67 117 69
rect 113 62 117 67
rect 113 60 114 62
rect 116 60 117 62
rect 73 48 75 49
rect 65 47 75 48
rect 77 47 78 49
rect 65 45 78 47
rect 65 43 67 45
rect 69 43 78 45
rect 65 42 78 43
rect 113 39 117 60
rect 93 38 117 39
rect 93 36 95 38
rect 97 36 117 38
rect 93 35 117 36
rect 121 71 126 73
rect 121 69 123 71
rect 125 69 126 71
rect 161 74 173 80
rect 121 64 126 69
rect 121 62 123 64
rect 125 62 126 64
rect 121 60 126 62
rect 153 69 157 72
rect 153 67 154 69
rect 156 67 157 69
rect 121 54 125 60
rect 121 52 122 54
rect 124 52 125 54
rect 121 40 125 52
rect 153 63 157 67
rect 144 62 157 63
rect 144 60 145 62
rect 147 60 150 62
rect 152 60 157 62
rect 144 59 157 60
rect 161 69 166 74
rect 161 67 163 69
rect 165 67 166 69
rect 161 62 166 67
rect 161 60 163 62
rect 165 60 166 62
rect 161 58 166 60
rect 136 54 150 55
rect 136 52 140 54
rect 142 52 150 54
rect 136 51 150 52
rect 121 38 123 40
rect 125 38 133 40
rect 121 34 133 38
rect 145 45 150 51
rect 145 43 146 45
rect 148 43 150 45
rect 145 42 150 43
rect 177 49 182 56
rect 205 71 221 72
rect 205 69 207 71
rect 209 69 221 71
rect 205 67 221 69
rect 177 48 179 49
rect 169 47 179 48
rect 181 47 182 49
rect 169 45 182 47
rect 169 43 171 45
rect 173 43 182 45
rect 169 42 182 43
rect 217 50 221 67
rect 234 63 238 72
rect 314 79 318 80
rect 305 75 318 79
rect 265 71 270 73
rect 234 62 247 63
rect 234 60 239 62
rect 241 60 247 62
rect 234 59 247 60
rect 217 48 218 50
rect 220 48 221 50
rect 217 39 221 48
rect 241 54 255 55
rect 241 52 249 54
rect 251 52 255 54
rect 241 51 255 52
rect 265 69 266 71
rect 268 69 270 71
rect 265 64 270 69
rect 265 62 266 64
rect 268 62 270 64
rect 265 60 270 62
rect 241 42 246 51
rect 266 59 270 60
rect 282 63 286 72
rect 282 61 303 63
rect 282 59 287 61
rect 289 59 303 61
rect 266 57 267 59
rect 269 57 270 59
rect 266 40 270 57
rect 282 54 303 55
rect 282 52 297 54
rect 299 52 303 54
rect 282 51 303 52
rect 316 73 318 75
rect 314 68 318 73
rect 316 66 318 68
rect 282 42 286 51
rect 314 60 318 66
rect 314 58 315 60
rect 317 58 318 60
rect 314 47 318 58
rect 313 45 318 47
rect 313 43 314 45
rect 316 43 318 45
rect 313 41 318 43
rect 331 78 344 79
rect 331 76 333 78
rect 335 76 344 78
rect 331 75 344 76
rect 331 52 335 75
rect 386 74 391 80
rect 386 72 387 74
rect 389 72 391 74
rect 331 50 332 52
rect 334 50 335 52
rect 386 71 391 72
rect 378 67 391 71
rect 405 78 418 79
rect 405 76 407 78
rect 409 76 418 78
rect 405 75 418 76
rect 340 56 342 58
rect 331 42 335 50
rect 346 62 359 64
rect 346 60 347 62
rect 349 60 359 62
rect 346 59 359 60
rect 346 57 347 59
rect 349 58 359 59
rect 376 61 378 63
rect 349 57 351 58
rect 346 50 351 57
rect 371 52 378 56
rect 371 50 374 52
rect 376 50 378 52
rect 371 49 378 50
rect 371 47 374 49
rect 376 47 378 49
rect 371 43 384 47
rect 197 38 221 39
rect 197 36 199 38
rect 201 36 221 38
rect 197 35 221 36
rect 258 38 266 40
rect 268 38 270 40
rect 258 34 270 38
rect 331 40 336 42
rect 331 38 333 40
rect 335 38 336 40
rect 331 36 336 38
rect 331 34 335 36
rect 405 56 409 75
rect 460 74 465 80
rect 460 72 461 74
rect 463 72 465 74
rect 405 54 406 56
rect 408 54 409 56
rect 405 42 409 54
rect 460 71 465 72
rect 452 67 465 71
rect 479 78 492 79
rect 479 76 481 78
rect 483 76 492 78
rect 479 75 492 76
rect 421 61 433 64
rect 414 56 416 58
rect 420 59 433 61
rect 420 57 421 59
rect 423 58 433 59
rect 450 61 452 63
rect 423 57 427 58
rect 420 55 427 57
rect 421 54 427 55
rect 421 52 423 54
rect 425 52 427 54
rect 421 50 427 52
rect 445 54 451 56
rect 445 52 448 54
rect 450 52 451 54
rect 445 47 451 52
rect 445 43 458 47
rect 405 40 410 42
rect 405 38 407 40
rect 409 38 410 40
rect 405 36 410 38
rect 405 34 409 36
rect 479 42 483 75
rect 534 74 539 80
rect 534 72 535 74
rect 537 72 539 74
rect 534 71 539 72
rect 526 67 539 71
rect 488 56 490 58
rect 495 59 507 64
rect 497 58 507 59
rect 524 61 526 63
rect 497 57 499 58
rect 495 56 499 57
rect 495 54 496 56
rect 498 54 499 56
rect 495 50 499 54
rect 519 54 525 56
rect 519 52 522 54
rect 524 52 525 54
rect 519 47 525 52
rect 519 45 522 47
rect 524 45 532 47
rect 519 43 532 45
rect 479 40 484 42
rect 479 38 481 40
rect 483 38 484 40
rect 479 36 484 38
rect 479 34 483 36
rect -27 28 543 29
rect -27 26 -20 28
rect -18 26 20 28
rect 22 26 30 28
rect 32 26 60 28
rect 62 26 113 28
rect 115 26 124 28
rect 126 26 134 28
rect 136 26 164 28
rect 166 26 217 28
rect 219 26 255 28
rect 257 26 265 28
rect 267 26 313 28
rect 315 26 543 28
rect -27 21 543 26
<< alu2 >>
rect 399 87 525 91
rect 226 80 393 84
rect 49 69 62 70
rect 9 67 22 69
rect 9 65 10 67
rect 12 65 18 67
rect 20 65 22 67
rect 49 67 50 69
rect 52 67 59 69
rect 61 67 62 69
rect 49 66 62 67
rect 153 69 166 70
rect 153 67 154 69
rect 156 67 163 69
rect 165 67 166 69
rect 153 66 166 67
rect 9 64 22 65
rect 113 62 148 63
rect 113 60 114 62
rect 116 60 145 62
rect 147 60 148 62
rect 113 59 148 60
rect 9 54 125 55
rect 9 52 10 54
rect 12 52 122 54
rect 124 52 125 54
rect 9 51 125 52
rect 226 51 230 80
rect 270 68 377 72
rect 270 60 275 68
rect 346 62 351 64
rect 346 61 347 62
rect 266 59 275 60
rect 266 57 267 59
rect 269 57 275 59
rect 314 60 347 61
rect 349 60 351 62
rect 314 58 315 60
rect 317 58 351 60
rect 314 57 351 58
rect 266 56 275 57
rect 346 56 350 57
rect 217 50 230 51
rect 217 48 218 50
rect 220 48 230 50
rect 217 47 230 48
rect 327 52 335 53
rect 327 50 332 52
rect 334 50 335 52
rect 327 49 335 50
rect 373 52 377 68
rect 373 50 374 52
rect 376 50 377 52
rect 41 45 73 47
rect 41 43 42 45
rect 44 43 67 45
rect 69 43 73 45
rect 41 42 73 43
rect 145 45 177 47
rect 145 43 146 45
rect 148 43 171 45
rect 173 43 177 45
rect 145 42 177 43
rect 327 27 331 49
rect 373 47 377 50
rect 389 38 393 80
rect 399 57 403 87
rect 399 56 409 57
rect 399 54 406 56
rect 408 54 409 56
rect 399 53 409 54
rect 422 54 426 60
rect 422 52 423 54
rect 425 52 426 54
rect 422 38 426 52
rect 389 34 426 38
rect 495 56 499 61
rect 495 54 496 56
rect 498 54 499 56
rect 495 27 499 54
rect 521 47 525 87
rect 521 45 522 47
rect 524 45 525 47
rect 521 44 525 45
rect 327 23 499 27
<< ptie >>
rect -22 28 -16 30
rect 18 28 24 30
rect -22 26 -20 28
rect -18 26 -16 28
rect -22 24 -16 26
rect 18 26 20 28
rect 22 26 24 28
rect 18 24 24 26
rect 58 28 64 30
rect 58 26 60 28
rect 62 26 64 28
rect 58 24 64 26
rect 122 28 128 30
rect 122 26 124 28
rect 126 26 128 28
rect 122 24 128 26
rect 162 28 168 30
rect 162 26 164 28
rect 166 26 168 28
rect 162 24 168 26
rect 263 28 269 30
rect 311 28 317 30
rect 263 26 265 28
rect 267 26 269 28
rect 263 24 269 26
rect 311 26 313 28
rect 315 26 317 28
rect 311 24 317 26
<< ntie >>
rect -22 88 -16 90
rect -22 86 -20 88
rect -18 86 -16 88
rect 18 88 24 90
rect -22 84 -16 86
rect 18 86 20 88
rect 22 86 24 88
rect 91 88 97 90
rect 18 84 24 86
rect 91 86 93 88
rect 95 86 97 88
rect 122 88 128 90
rect 91 84 97 86
rect 122 86 124 88
rect 126 86 128 88
rect 195 88 201 90
rect 122 84 128 86
rect 195 86 197 88
rect 199 86 201 88
rect 263 88 269 90
rect 195 84 201 86
rect 263 86 265 88
rect 267 86 269 88
rect 311 88 317 90
rect 263 84 269 86
rect 311 86 313 88
rect 315 86 317 88
rect 311 84 317 86
<< nmos >>
rect -16 38 -14 47
rect -6 41 -4 47
rect 4 41 6 47
rect 24 36 26 45
rect 37 34 39 45
rect 44 34 46 45
rect 64 38 66 47
rect 80 33 82 42
rect 90 33 92 42
rect 100 30 102 42
rect 107 30 109 42
rect 128 36 130 45
rect 141 34 143 45
rect 148 34 150 45
rect 168 38 170 47
rect 184 33 186 42
rect 194 33 196 42
rect 204 30 206 42
rect 211 30 213 42
rect 241 34 243 45
rect 248 34 250 45
rect 261 36 263 45
rect 289 41 291 47
rect 299 41 301 47
rect 309 38 311 47
rect 338 33 340 42
rect 348 33 350 41
rect 355 33 357 41
rect 365 33 367 41
rect 372 33 374 41
rect 382 35 384 41
rect 412 33 414 42
rect 422 33 424 41
rect 429 33 431 41
rect 439 33 441 41
rect 446 33 448 41
rect 456 35 458 41
rect 486 33 488 42
rect 496 33 498 41
rect 503 33 505 41
rect 513 33 515 41
rect 520 33 522 41
rect 530 35 532 41
<< pmos >>
rect -16 59 -14 77
rect -3 66 -1 87
rect 4 66 6 87
rect 24 60 26 78
rect 34 67 36 80
rect 44 67 46 80
rect 72 60 74 87
rect 88 60 90 78
rect 98 60 100 78
rect 108 60 110 87
rect 128 60 130 78
rect 138 67 140 80
rect 148 67 150 80
rect 176 60 178 87
rect 192 60 194 78
rect 202 60 204 78
rect 212 60 214 87
rect 241 67 243 80
rect 251 67 253 80
rect 261 60 263 78
rect 289 66 291 87
rect 296 66 298 87
rect 309 59 311 77
rect 338 69 340 87
rect 348 71 350 87
rect 355 71 357 87
rect 365 71 367 87
rect 372 71 374 87
rect 412 69 414 87
rect 422 71 424 87
rect 429 71 431 87
rect 439 71 441 87
rect 446 71 448 87
rect 382 59 384 67
rect 486 69 488 87
rect 496 71 498 87
rect 503 71 505 87
rect 513 71 515 87
rect 520 71 522 87
rect 456 59 458 67
rect 530 59 532 67
<< polyct0 >>
rect -14 52 -12 54
rect 26 52 28 54
rect 96 52 98 54
rect 106 53 108 55
rect 130 52 132 54
rect 200 52 202 54
rect 210 53 212 55
rect 259 52 261 54
rect 307 52 309 54
rect 364 62 366 64
rect 339 47 341 49
rect 357 46 359 48
rect 438 62 440 64
rect 413 47 415 49
rect 431 46 433 48
rect 512 62 514 64
rect 487 47 489 49
rect 505 46 507 48
<< polyct1 >>
rect 6 59 8 61
rect -4 52 -2 54
rect 46 60 48 62
rect 59 60 61 62
rect 36 52 38 54
rect 150 60 152 62
rect 163 60 165 62
rect 239 60 241 62
rect 75 47 77 49
rect 140 52 142 54
rect 179 47 181 49
rect 287 59 289 61
rect 249 52 251 54
rect 387 72 389 74
rect 297 52 299 54
rect 347 57 349 59
rect 461 72 463 74
rect 374 47 376 49
rect 421 57 423 59
rect 535 72 537 74
rect 448 52 450 54
rect 495 57 497 59
rect 522 52 524 54
<< ndifct0 >>
rect -1 43 1 45
rect -10 30 -8 32
rect 59 43 61 45
rect 49 36 51 38
rect 73 35 75 37
rect 9 30 11 32
rect 85 38 87 40
rect 163 43 165 45
rect 153 36 155 38
rect 177 35 179 37
rect 189 38 191 40
rect 236 36 238 38
rect 294 43 296 45
rect 284 30 286 32
rect 343 35 345 37
rect 360 35 362 37
rect 377 37 379 39
rect 387 37 389 39
rect 303 30 305 32
rect 417 35 419 37
rect 434 35 436 37
rect 451 37 453 39
rect 461 37 463 39
rect 491 35 493 37
rect 508 35 510 37
rect 525 37 527 39
rect 535 37 537 39
<< ndifct1 >>
rect -21 43 -19 45
rect 19 38 21 40
rect 95 36 97 38
rect 30 26 32 28
rect 123 38 125 40
rect 113 26 115 28
rect 199 36 201 38
rect 134 26 136 28
rect 266 38 268 40
rect 217 26 219 28
rect 314 43 316 45
rect 333 38 335 40
rect 255 26 257 28
rect 407 38 409 40
rect 481 38 483 40
<< ntiect1 >>
rect -20 86 -18 88
rect 20 86 22 88
rect 93 86 95 88
rect 124 86 126 88
rect 197 86 199 88
rect 265 86 267 88
rect 313 86 315 88
<< ptiect1 >>
rect -20 26 -18 28
rect 20 26 22 28
rect 60 26 62 28
rect 124 26 126 28
rect 164 26 166 28
rect 265 26 267 28
rect 313 26 315 28
<< pdifct0 >>
rect -10 83 -8 85
rect 9 76 11 78
rect 29 74 31 76
rect 39 76 41 78
rect 39 69 41 71
rect 49 76 51 78
rect 67 62 69 64
rect 77 83 79 85
rect 77 76 79 78
rect 93 69 95 71
rect 93 62 95 64
rect 113 77 115 79
rect 133 74 135 76
rect 143 76 145 78
rect 143 69 145 71
rect 153 76 155 78
rect 171 62 173 64
rect 181 83 183 85
rect 181 76 183 78
rect 197 69 199 71
rect 197 62 199 64
rect 217 77 219 79
rect 236 76 238 78
rect 246 76 248 78
rect 246 69 248 71
rect 256 74 258 76
rect 284 76 286 78
rect 303 83 305 85
rect 343 83 345 85
rect 360 73 362 75
rect 377 83 379 85
rect 417 83 419 85
rect 434 73 436 75
rect 451 83 453 85
rect 387 61 389 63
rect 491 83 493 85
rect 508 73 510 75
rect 525 83 527 85
rect 461 61 463 63
rect 535 61 537 63
<< pdifct1 >>
rect -21 73 -19 75
rect -21 66 -19 68
rect 19 69 21 71
rect 19 62 21 64
rect 103 69 105 71
rect 123 69 125 71
rect 123 62 125 64
rect 207 69 209 71
rect 266 69 268 71
rect 266 62 268 64
rect 314 73 316 75
rect 333 76 335 78
rect 407 76 409 78
rect 314 66 316 68
rect 481 76 483 78
<< alu0 >>
rect -12 83 -10 85
rect -8 83 -6 85
rect -12 82 -6 83
rect -4 78 13 79
rect -4 76 9 78
rect 11 76 13 78
rect -4 75 13 76
rect 27 76 33 85
rect -19 64 -18 75
rect -4 71 0 75
rect 27 74 29 76
rect 31 74 33 76
rect 27 73 33 74
rect 38 78 42 80
rect 38 76 39 78
rect 41 76 42 78
rect -15 67 0 71
rect -15 54 -11 67
rect 38 71 42 76
rect 47 78 53 85
rect 76 83 77 85
rect 79 83 80 85
rect 47 76 49 78
rect 51 76 53 78
rect 47 75 53 76
rect 76 78 80 83
rect 76 76 77 78
rect 79 76 80 78
rect 76 74 80 76
rect 84 79 117 80
rect 84 77 113 79
rect 115 77 117 79
rect 84 76 117 77
rect 131 76 137 85
rect 38 70 39 71
rect 25 69 39 70
rect 41 69 42 71
rect 25 66 42 69
rect 4 58 10 59
rect -15 52 -14 54
rect -12 52 -11 54
rect -15 46 -11 52
rect -15 45 3 46
rect -15 43 -1 45
rect 1 43 3 45
rect -15 42 3 43
rect 25 54 29 66
rect 84 65 88 76
rect 131 74 133 76
rect 135 74 137 76
rect 131 73 137 74
rect 142 78 146 80
rect 142 76 143 78
rect 145 76 146 78
rect 65 64 88 65
rect 65 62 67 64
rect 69 62 88 64
rect 65 61 88 62
rect 65 55 69 61
rect 25 52 26 54
rect 28 52 29 54
rect 25 47 29 52
rect 25 43 37 47
rect 21 40 22 42
rect 33 39 37 43
rect 58 51 69 55
rect 58 45 62 51
rect 84 55 88 61
rect 92 71 96 73
rect 92 69 93 71
rect 95 69 96 71
rect 92 64 96 69
rect 92 62 93 64
rect 95 63 96 64
rect 95 62 108 63
rect 92 59 108 62
rect 104 57 108 59
rect 104 55 109 57
rect 84 54 100 55
rect 84 52 96 54
rect 98 52 100 54
rect 84 51 100 52
rect 104 53 106 55
rect 108 53 109 55
rect 104 51 109 53
rect 58 43 59 45
rect 61 43 62 45
rect 58 41 62 43
rect 104 47 108 51
rect 84 43 108 47
rect 84 40 88 43
rect 33 38 53 39
rect 84 38 85 40
rect 87 38 88 40
rect 33 36 49 38
rect 51 36 53 38
rect 33 35 53 36
rect 71 37 77 38
rect 71 35 73 37
rect 75 35 77 37
rect 84 36 88 38
rect 142 71 146 76
rect 151 78 157 85
rect 180 83 181 85
rect 183 83 184 85
rect 151 76 153 78
rect 155 76 157 78
rect 151 75 157 76
rect 180 78 184 83
rect 180 76 181 78
rect 183 76 184 78
rect 180 74 184 76
rect 188 79 221 80
rect 188 77 217 79
rect 219 77 221 79
rect 188 76 221 77
rect 234 78 240 85
rect 234 76 236 78
rect 238 76 240 78
rect 142 70 143 71
rect 129 69 143 70
rect 145 69 146 71
rect 129 66 146 69
rect 129 54 133 66
rect 188 65 192 76
rect 234 75 240 76
rect 245 78 249 80
rect 245 76 246 78
rect 248 76 249 78
rect 169 64 192 65
rect 169 62 171 64
rect 173 62 192 64
rect 169 61 192 62
rect 169 55 173 61
rect 129 52 130 54
rect 132 52 133 54
rect 129 47 133 52
rect 129 43 141 47
rect 125 40 126 42
rect -12 32 -6 33
rect -12 30 -10 32
rect -8 30 -6 32
rect -12 29 -6 30
rect 7 32 13 33
rect 7 30 9 32
rect 11 30 13 32
rect 7 29 13 30
rect 71 29 77 35
rect 137 39 141 43
rect 162 51 173 55
rect 162 45 166 51
rect 188 55 192 61
rect 196 71 200 73
rect 196 69 197 71
rect 199 69 200 71
rect 196 64 200 69
rect 196 62 197 64
rect 199 63 200 64
rect 199 62 212 63
rect 196 59 212 62
rect 208 57 212 59
rect 208 55 213 57
rect 188 54 204 55
rect 188 52 200 54
rect 202 52 204 54
rect 188 51 204 52
rect 208 53 210 55
rect 212 53 213 55
rect 208 51 213 53
rect 162 43 163 45
rect 165 43 166 45
rect 162 41 166 43
rect 208 47 212 51
rect 188 43 212 47
rect 245 71 249 76
rect 254 76 260 85
rect 301 83 303 85
rect 305 83 307 85
rect 301 82 307 83
rect 341 83 343 85
rect 345 83 347 85
rect 341 82 347 83
rect 376 83 377 85
rect 379 83 380 85
rect 376 81 380 83
rect 415 83 417 85
rect 419 83 421 85
rect 415 82 421 83
rect 450 83 451 85
rect 453 83 454 85
rect 450 81 454 83
rect 489 83 491 85
rect 493 83 495 85
rect 489 82 495 83
rect 524 83 525 85
rect 527 83 528 85
rect 524 81 528 83
rect 254 74 256 76
rect 258 74 260 76
rect 282 78 299 79
rect 282 76 284 78
rect 286 76 299 78
rect 282 75 299 76
rect 254 73 260 74
rect 245 69 246 71
rect 248 70 249 71
rect 248 69 262 70
rect 245 66 262 69
rect 188 40 192 43
rect 137 38 157 39
rect 188 38 189 40
rect 191 38 192 40
rect 258 54 262 66
rect 258 52 259 54
rect 261 52 262 54
rect 258 47 262 52
rect 250 43 262 47
rect 295 71 299 75
rect 295 67 310 71
rect 285 58 291 59
rect 250 39 254 43
rect 265 40 266 42
rect 306 54 310 67
rect 313 64 314 75
rect 306 52 307 54
rect 309 52 310 54
rect 306 46 310 52
rect 292 45 310 46
rect 292 43 294 45
rect 296 43 310 45
rect 292 42 310 43
rect 351 75 364 76
rect 351 73 360 75
rect 362 73 364 75
rect 351 72 364 73
rect 339 68 355 72
rect 339 58 343 68
rect 425 75 438 76
rect 363 64 367 66
rect 339 56 340 58
rect 342 56 343 58
rect 339 51 343 56
rect 338 49 343 51
rect 363 62 364 64
rect 366 63 391 64
rect 366 62 376 63
rect 363 61 376 62
rect 378 61 387 63
rect 389 61 391 63
rect 363 60 391 61
rect 363 50 367 60
rect 338 47 339 49
rect 341 47 343 49
rect 356 48 367 50
rect 338 45 353 47
rect 339 43 353 45
rect 356 46 357 48
rect 359 46 367 48
rect 356 44 367 46
rect 137 36 153 38
rect 155 36 157 38
rect 137 35 157 36
rect 175 37 181 38
rect 175 35 177 37
rect 179 35 181 37
rect 188 36 192 38
rect 234 38 254 39
rect 234 36 236 38
rect 238 36 254 38
rect 234 35 254 36
rect 175 29 181 35
rect 342 37 346 39
rect 342 35 343 37
rect 345 35 346 37
rect 282 32 288 33
rect 282 30 284 32
rect 286 30 288 32
rect 282 29 288 30
rect 301 32 307 33
rect 301 30 303 32
rect 305 30 307 32
rect 301 29 307 30
rect 342 29 346 35
rect 349 38 353 43
rect 387 40 391 60
rect 375 39 381 40
rect 349 37 364 38
rect 349 35 360 37
rect 362 35 364 37
rect 349 34 364 35
rect 375 37 377 39
rect 379 37 381 39
rect 375 29 381 37
rect 385 39 391 40
rect 385 37 387 39
rect 389 37 391 39
rect 385 36 391 37
rect 425 73 434 75
rect 436 73 438 75
rect 425 72 438 73
rect 413 68 429 72
rect 413 58 417 68
rect 499 75 512 76
rect 437 64 441 66
rect 413 56 414 58
rect 416 56 417 58
rect 413 51 417 56
rect 437 62 438 64
rect 440 63 465 64
rect 440 62 450 63
rect 437 61 450 62
rect 452 61 461 63
rect 463 61 465 63
rect 437 60 465 61
rect 412 49 417 51
rect 437 50 441 60
rect 412 47 413 49
rect 415 47 417 49
rect 430 48 441 50
rect 412 45 427 47
rect 413 43 427 45
rect 430 46 431 48
rect 433 46 441 48
rect 430 44 441 46
rect 416 37 420 39
rect 416 35 417 37
rect 419 35 420 37
rect 416 29 420 35
rect 423 38 427 43
rect 461 40 465 60
rect 449 39 455 40
rect 423 37 438 38
rect 423 35 434 37
rect 436 35 438 37
rect 423 34 438 35
rect 449 37 451 39
rect 453 37 455 39
rect 449 29 455 37
rect 459 39 465 40
rect 459 37 461 39
rect 463 37 465 39
rect 459 36 465 37
rect 499 73 508 75
rect 510 73 512 75
rect 499 72 512 73
rect 487 68 503 72
rect 487 58 491 68
rect 511 64 515 66
rect 487 56 488 58
rect 490 56 491 58
rect 487 51 491 56
rect 494 55 495 61
rect 511 62 512 64
rect 514 63 539 64
rect 514 62 524 63
rect 511 61 524 62
rect 526 61 535 63
rect 537 61 539 63
rect 511 60 539 61
rect 486 49 491 51
rect 511 50 515 60
rect 486 47 487 49
rect 489 47 491 49
rect 504 48 515 50
rect 486 45 501 47
rect 487 43 501 45
rect 504 46 505 48
rect 507 46 515 48
rect 504 44 515 46
rect 490 37 494 39
rect 490 35 491 37
rect 493 35 494 37
rect 490 29 494 35
rect 497 38 501 43
rect 535 40 539 60
rect 523 39 529 40
rect 497 37 512 38
rect 497 35 508 37
rect 510 35 512 37
rect 497 34 512 35
rect 523 37 525 39
rect 527 37 529 39
rect 523 29 529 37
rect 533 39 539 40
rect 533 37 535 39
rect 537 37 539 39
rect 533 36 539 37
<< via1 >>
rect 10 65 12 67
rect 18 65 20 67
rect 50 67 52 69
rect 10 52 12 54
rect 59 67 61 69
rect 42 43 44 45
rect 114 60 116 62
rect 67 43 69 45
rect 154 67 156 69
rect 122 52 124 54
rect 145 60 147 62
rect 163 67 165 69
rect 146 43 148 45
rect 171 43 173 45
rect 218 48 220 50
rect 267 57 269 59
rect 315 58 317 60
rect 332 50 334 52
rect 347 60 349 62
rect 374 50 376 52
rect 406 54 408 56
rect 423 52 425 54
rect 496 54 498 56
rect 522 45 524 47
<< labels >>
rlabel alu0 60 48 60 48 6 bn
rlabel alu0 106 53 106 53 6 an
rlabel alu1 75 49 75 49 6 a
rlabel alu1 51 69 51 69 6 b
rlabel alu1 35 53 35 53 6 a
rlabel alu0 27 56 27 56 6 zn
rlabel via1 219 49 219 49 1 sum
rlabel alu1 115 49 115 49 1 s
rlabel alu1 139 52 139 52 1 cin
rlabel alu1 27 37 27 37 1 co
rlabel alu0 131 55 131 55 1 zn_1
rlabel alu0 164 48 164 48 1 bn_1
rlabel alu0 190 40 190 40 1 an_1
rlabel alu1 131 37 131 37 1 c1
rlabel alu1 -21 57 -21 57 1 cout
rlabel alu0 4 77 4 77 1 zn_2
rlabel polyct1 348 58 348 58 1 i0
rlabel polyct1 422 58 422 58 1 i2
rlabel polyct1 449 53 449 53 1 i3
rlabel polyct1 388 73 388 73 1 s0
rlabel polyct1 462 73 462 73 1 s0
rlabel polyct1 536 73 536 73 1 s1
rlabel alu1 389 90 389 90 1 vdd!
rlabel alu1 507 24 507 24 1 vss!
rlabel alu1 252 53 252 53 4 a
rlabel alu1 244 49 244 49 4 a
rlabel alu1 244 61 244 61 4 b
rlabel alu1 236 69 236 69 4 b
rlabel alu1 300 53 300 53 4 a
rlabel alu1 292 53 292 53 4 a
rlabel alu1 292 61 292 61 4 b
rlabel alu1 300 61 300 61 4 b
rlabel alu1 284 45 284 45 4 a
rlabel alu1 284 69 284 69 4 b
rlabel alu2 375 48 375 48 1 i1
rlabel alu1 481 56 481 56 1 aluout
<< end >>
