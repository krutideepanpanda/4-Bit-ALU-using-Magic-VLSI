magic
tech scmos
timestamp 1607366742
<< ab >>
rect -35 69 213 77
rect -35 37 45 69
rect 46 37 149 69
rect 150 37 213 69
rect -35 5 213 37
rect 40 0 46 5
rect 144 0 150 5
<< nwell >>
rect -40 37 218 82
<< pwell >>
rect -40 0 218 37
<< poly >>
rect -13 71 -11 75
rect -6 71 -4 75
rect -26 61 -24 66
rect 62 71 64 75
rect 14 62 16 66
rect 24 64 26 69
rect 34 64 36 69
rect -26 40 -24 43
rect -13 40 -11 50
rect -6 47 -4 50
rect -6 45 0 47
rect -6 43 -4 45
rect -2 43 0 45
rect -6 41 0 43
rect -26 38 -20 40
rect -26 36 -24 38
rect -22 36 -20 38
rect -26 34 -20 36
rect -16 38 -10 40
rect -16 36 -14 38
rect -12 36 -10 38
rect -16 34 -10 36
rect -26 31 -24 34
rect -16 31 -14 34
rect -6 31 -4 41
rect 14 40 16 44
rect 24 40 26 51
rect 34 48 36 51
rect 34 46 40 48
rect 34 44 36 46
rect 38 44 40 46
rect 34 42 40 44
rect 47 46 53 48
rect 47 44 49 46
rect 51 44 53 46
rect 98 71 100 75
rect 78 62 80 66
rect 88 62 90 66
rect 166 71 168 75
rect 118 62 120 66
rect 128 64 130 69
rect 138 64 140 69
rect 47 42 53 44
rect 14 38 20 40
rect 14 36 16 38
rect 18 36 20 38
rect 14 34 20 36
rect 24 38 30 40
rect 24 36 26 38
rect 28 36 30 38
rect 24 34 30 36
rect 14 29 16 34
rect 27 29 29 34
rect 34 29 36 42
rect 51 41 53 42
rect 62 41 64 44
rect 78 41 80 44
rect 51 39 64 41
rect 70 39 80 41
rect 88 40 90 44
rect 98 41 100 44
rect 54 31 56 39
rect 70 35 72 39
rect 63 33 72 35
rect 84 38 90 40
rect 84 36 86 38
rect 88 36 90 38
rect 84 34 90 36
rect 94 39 100 41
rect 94 37 96 39
rect 98 37 100 39
rect 94 35 100 37
rect 118 40 120 44
rect 128 40 130 51
rect 138 48 140 51
rect 138 46 144 48
rect 138 44 140 46
rect 142 44 144 46
rect 138 42 144 44
rect 151 46 157 48
rect 151 44 153 46
rect 155 44 157 46
rect 202 71 204 75
rect 182 62 184 66
rect 192 62 194 66
rect 151 42 157 44
rect 118 38 124 40
rect 118 36 120 38
rect 122 36 124 38
rect 63 31 65 33
rect 67 31 72 33
rect -26 17 -24 22
rect -16 20 -14 25
rect -6 20 -4 25
rect 14 16 16 20
rect 63 29 72 31
rect 88 31 90 34
rect 70 26 72 29
rect 80 26 82 30
rect 88 29 92 31
rect 90 26 92 29
rect 97 26 99 35
rect 118 34 124 36
rect 128 38 134 40
rect 128 36 130 38
rect 132 36 134 38
rect 128 34 134 36
rect 118 29 120 34
rect 131 29 133 34
rect 138 29 140 42
rect 155 41 157 42
rect 166 41 168 44
rect 182 41 184 44
rect 155 39 168 41
rect 174 39 184 41
rect 192 40 194 44
rect 202 41 204 44
rect 158 31 160 39
rect 174 35 176 39
rect 167 33 176 35
rect 188 38 194 40
rect 188 36 190 38
rect 192 36 194 38
rect 188 34 194 36
rect 198 39 204 41
rect 198 37 200 39
rect 202 37 204 39
rect 198 35 204 37
rect 167 31 169 33
rect 171 31 176 33
rect 54 19 56 22
rect 27 13 29 18
rect 34 13 36 18
rect 54 17 59 19
rect 57 9 59 17
rect 70 13 72 17
rect 80 9 82 17
rect 118 16 120 20
rect 167 29 176 31
rect 192 31 194 34
rect 174 26 176 29
rect 184 26 186 30
rect 192 29 196 31
rect 194 26 196 29
rect 201 26 203 35
rect 158 19 160 22
rect 90 9 92 14
rect 97 9 99 14
rect 57 7 82 9
rect 131 13 133 18
rect 138 13 140 18
rect 158 17 163 19
rect 161 9 163 17
rect 174 13 176 17
rect 184 9 186 17
rect 194 9 196 14
rect 201 9 203 14
rect 161 7 186 9
<< ndif >>
rect -33 29 -26 31
rect -33 27 -31 29
rect -29 27 -26 29
rect -33 25 -26 27
rect -31 22 -26 25
rect -24 25 -16 31
rect -14 29 -6 31
rect -14 27 -11 29
rect -9 27 -6 29
rect -14 25 -6 27
rect -4 25 3 31
rect 47 29 54 31
rect 9 26 14 29
rect -24 22 -18 25
rect -22 18 -18 22
rect -2 18 3 25
rect 7 24 14 26
rect 7 22 9 24
rect 11 22 14 24
rect 7 20 14 22
rect 16 20 27 29
rect -22 16 -16 18
rect -22 14 -20 16
rect -18 14 -16 16
rect -22 12 -16 14
rect -3 16 3 18
rect 18 18 27 20
rect 29 18 34 29
rect 36 24 41 29
rect 47 27 49 29
rect 51 27 54 29
rect 47 25 54 27
rect 36 22 43 24
rect 49 22 54 25
rect 56 26 61 31
rect 151 29 158 31
rect 113 26 118 29
rect 56 22 70 26
rect 36 20 39 22
rect 41 20 43 22
rect 36 18 43 20
rect 61 21 70 22
rect 61 19 63 21
rect 65 19 70 21
rect -3 14 -1 16
rect 1 14 3 16
rect -3 12 3 14
rect 18 12 25 18
rect 61 17 70 19
rect 72 24 80 26
rect 72 22 75 24
rect 77 22 80 24
rect 72 17 80 22
rect 82 22 90 26
rect 82 20 85 22
rect 87 20 90 22
rect 82 17 90 20
rect 18 10 20 12
rect 22 10 25 12
rect 18 8 25 10
rect 85 14 90 17
rect 92 14 97 26
rect 99 14 107 26
rect 111 24 118 26
rect 111 22 113 24
rect 115 22 118 24
rect 111 20 118 22
rect 120 20 131 29
rect 122 18 131 20
rect 133 18 138 29
rect 140 24 145 29
rect 151 27 153 29
rect 155 27 158 29
rect 151 25 158 27
rect 140 22 147 24
rect 153 22 158 25
rect 160 26 165 31
rect 160 22 174 26
rect 140 20 143 22
rect 145 20 147 22
rect 140 18 147 20
rect 165 21 174 22
rect 165 19 167 21
rect 169 19 174 21
rect 101 12 107 14
rect 101 10 103 12
rect 105 10 107 12
rect 101 8 107 10
rect 122 12 129 18
rect 165 17 174 19
rect 176 24 184 26
rect 176 22 179 24
rect 181 22 184 24
rect 176 17 184 22
rect 186 22 194 26
rect 186 20 189 22
rect 191 20 194 22
rect 186 17 194 20
rect 122 10 124 12
rect 126 10 129 12
rect 122 8 129 10
rect 189 14 194 17
rect 196 14 201 26
rect 203 14 211 26
rect 205 12 211 14
rect 205 10 207 12
rect 209 10 211 12
rect 205 8 211 10
<< pdif >>
rect -22 69 -13 71
rect -22 67 -20 69
rect -18 67 -13 69
rect -22 61 -13 67
rect -33 59 -26 61
rect -33 57 -31 59
rect -29 57 -26 59
rect -33 52 -26 57
rect -33 50 -31 52
rect -29 50 -26 52
rect -33 48 -26 50
rect -31 43 -26 48
rect -24 50 -13 61
rect -11 50 -6 71
rect -4 64 1 71
rect -4 62 3 64
rect 18 62 24 64
rect -4 60 -1 62
rect 1 60 3 62
rect -4 58 3 60
rect -4 50 1 58
rect 9 57 14 62
rect 7 55 14 57
rect 7 53 9 55
rect 11 53 14 55
rect -24 43 -16 50
rect 7 48 14 53
rect 7 46 9 48
rect 11 46 14 48
rect 7 44 14 46
rect 16 60 24 62
rect 16 58 19 60
rect 21 58 24 60
rect 16 51 24 58
rect 26 62 34 64
rect 26 60 29 62
rect 31 60 34 62
rect 26 55 34 60
rect 26 53 29 55
rect 31 53 34 55
rect 26 51 34 53
rect 36 62 43 64
rect 36 60 39 62
rect 41 60 43 62
rect 36 51 43 60
rect 16 44 22 51
rect 57 50 62 71
rect 55 48 62 50
rect 55 46 57 48
rect 59 46 62 48
rect 55 44 62 46
rect 64 69 76 71
rect 64 67 67 69
rect 69 67 76 69
rect 64 62 76 67
rect 93 62 98 71
rect 64 60 67 62
rect 69 60 78 62
rect 64 44 78 60
rect 80 55 88 62
rect 80 53 83 55
rect 85 53 88 55
rect 80 48 88 53
rect 80 46 83 48
rect 85 46 88 48
rect 80 44 88 46
rect 90 55 98 62
rect 90 53 93 55
rect 95 53 98 55
rect 90 44 98 53
rect 100 65 105 71
rect 100 63 107 65
rect 100 61 103 63
rect 105 61 107 63
rect 122 62 128 64
rect 100 59 107 61
rect 100 44 105 59
rect 113 57 118 62
rect 111 55 118 57
rect 111 53 113 55
rect 115 53 118 55
rect 111 48 118 53
rect 111 46 113 48
rect 115 46 118 48
rect 111 44 118 46
rect 120 60 128 62
rect 120 58 123 60
rect 125 58 128 60
rect 120 51 128 58
rect 130 62 138 64
rect 130 60 133 62
rect 135 60 138 62
rect 130 55 138 60
rect 130 53 133 55
rect 135 53 138 55
rect 130 51 138 53
rect 140 62 147 64
rect 140 60 143 62
rect 145 60 147 62
rect 140 51 147 60
rect 120 44 126 51
rect 161 50 166 71
rect 159 48 166 50
rect 159 46 161 48
rect 163 46 166 48
rect 159 44 166 46
rect 168 69 180 71
rect 168 67 171 69
rect 173 67 180 69
rect 168 62 180 67
rect 197 62 202 71
rect 168 60 171 62
rect 173 60 182 62
rect 168 44 182 60
rect 184 55 192 62
rect 184 53 187 55
rect 189 53 192 55
rect 184 48 192 53
rect 184 46 187 48
rect 189 46 192 48
rect 184 44 192 46
rect 194 55 202 62
rect 194 53 197 55
rect 199 53 202 55
rect 194 44 202 53
rect 204 65 209 71
rect 204 63 211 65
rect 204 61 207 63
rect 209 61 211 63
rect 204 59 211 61
rect 204 44 209 59
<< alu1 >>
rect -37 72 215 77
rect -37 70 -30 72
rect -28 70 10 72
rect 12 70 83 72
rect 85 70 114 72
rect 116 70 187 72
rect 189 70 215 72
rect -37 69 215 70
rect -33 63 -29 64
rect -33 59 -20 63
rect -33 57 -31 59
rect -33 52 -29 57
rect -33 50 -31 52
rect -33 31 -29 50
rect -1 51 3 56
rect -1 49 0 51
rect 2 49 3 51
rect -1 47 3 49
rect -18 45 3 47
rect -18 43 -4 45
rect -2 43 3 45
rect 7 55 12 57
rect 7 53 9 55
rect 11 53 12 55
rect 47 58 59 64
rect 7 51 12 53
rect 7 49 8 51
rect 10 49 12 51
rect 7 48 12 49
rect 7 46 9 48
rect 11 46 12 48
rect 7 44 12 46
rect 39 53 43 56
rect 39 51 40 53
rect 42 51 43 53
rect -33 29 -28 31
rect -33 27 -31 29
rect -29 27 -28 29
rect -33 25 -28 27
rect -18 38 3 39
rect -18 36 -14 38
rect -12 36 0 38
rect 2 36 3 38
rect -18 35 3 36
rect -1 26 3 35
rect 7 24 11 44
rect 39 47 43 51
rect 30 46 43 47
rect 30 44 36 46
rect 38 44 43 46
rect 30 43 43 44
rect 47 53 52 58
rect 47 51 49 53
rect 51 51 52 53
rect 47 46 52 51
rect 47 44 49 46
rect 51 44 52 46
rect 47 42 52 44
rect 22 38 36 39
rect 22 36 26 38
rect 28 36 36 38
rect 22 35 36 36
rect 7 22 9 24
rect 11 22 19 24
rect 7 18 19 22
rect 31 29 36 35
rect 31 27 32 29
rect 34 27 36 29
rect 31 26 36 27
rect 63 33 68 40
rect 91 55 107 56
rect 91 53 93 55
rect 95 53 107 55
rect 91 51 107 53
rect 103 46 107 51
rect 103 44 104 46
rect 106 44 107 46
rect 63 32 65 33
rect 55 31 65 32
rect 67 31 68 33
rect 55 29 68 31
rect 55 27 57 29
rect 59 27 68 29
rect 55 26 68 27
rect 103 23 107 44
rect 83 22 107 23
rect 83 20 85 22
rect 87 20 107 22
rect 83 19 107 20
rect 111 55 116 57
rect 111 53 113 55
rect 115 53 116 55
rect 151 58 163 64
rect 111 48 116 53
rect 111 46 113 48
rect 115 46 116 48
rect 111 44 116 46
rect 143 53 147 56
rect 143 51 144 53
rect 146 51 147 53
rect 111 38 115 44
rect 111 36 112 38
rect 114 36 115 38
rect 111 24 115 36
rect 143 47 147 51
rect 134 46 147 47
rect 134 44 135 46
rect 137 44 140 46
rect 142 44 147 46
rect 134 43 147 44
rect 151 53 156 58
rect 151 51 153 53
rect 155 51 156 53
rect 151 46 156 51
rect 151 44 153 46
rect 155 44 156 46
rect 151 42 156 44
rect 126 38 140 39
rect 126 36 130 38
rect 132 36 140 38
rect 126 35 140 36
rect 111 22 113 24
rect 115 22 123 24
rect 111 18 123 22
rect 135 29 140 35
rect 135 27 136 29
rect 138 27 140 29
rect 135 26 140 27
rect 167 33 172 40
rect 195 55 211 56
rect 195 53 197 55
rect 199 53 211 55
rect 195 51 211 53
rect 167 32 169 33
rect 159 31 169 32
rect 171 31 172 33
rect 159 29 172 31
rect 159 27 161 29
rect 163 27 172 29
rect 159 26 172 27
rect 207 23 211 51
rect 187 22 211 23
rect 187 20 189 22
rect 191 20 211 22
rect 187 19 211 20
rect -37 12 215 13
rect -37 10 -30 12
rect -28 10 10 12
rect 12 10 20 12
rect 22 10 50 12
rect 52 10 103 12
rect 105 10 114 12
rect 116 10 124 12
rect 126 10 154 12
rect 156 10 207 12
rect 209 10 215 12
rect -37 5 215 10
<< alu2 >>
rect 39 53 52 54
rect -1 51 12 53
rect -1 49 0 51
rect 2 49 8 51
rect 10 49 12 51
rect 39 51 40 53
rect 42 51 49 53
rect 51 51 52 53
rect 39 50 52 51
rect 143 53 156 54
rect 143 51 144 53
rect 146 51 153 53
rect 155 51 156 53
rect 143 50 156 51
rect -1 48 12 49
rect 103 46 138 47
rect 103 44 104 46
rect 106 44 135 46
rect 137 44 138 46
rect 103 43 138 44
rect -1 38 115 39
rect -1 36 0 38
rect 2 36 112 38
rect 114 36 115 38
rect -1 35 115 36
rect 31 29 63 31
rect 31 27 32 29
rect 34 27 57 29
rect 59 27 63 29
rect 31 26 63 27
rect 135 29 167 31
rect 135 27 136 29
rect 138 27 161 29
rect 163 27 167 29
rect 135 26 167 27
<< ptie >>
rect -32 12 -26 14
rect 8 12 14 14
rect -32 10 -30 12
rect -28 10 -26 12
rect -32 8 -26 10
rect 8 10 10 12
rect 12 10 14 12
rect 8 8 14 10
rect 48 12 54 14
rect 48 10 50 12
rect 52 10 54 12
rect 48 8 54 10
rect 112 12 118 14
rect 112 10 114 12
rect 116 10 118 12
rect 112 8 118 10
rect 152 12 158 14
rect 152 10 154 12
rect 156 10 158 12
rect 152 8 158 10
<< ntie >>
rect -32 72 -26 74
rect -32 70 -30 72
rect -28 70 -26 72
rect 8 72 14 74
rect -32 68 -26 70
rect 8 70 10 72
rect 12 70 14 72
rect 81 72 87 74
rect 8 68 14 70
rect 81 70 83 72
rect 85 70 87 72
rect 112 72 118 74
rect 81 68 87 70
rect 112 70 114 72
rect 116 70 118 72
rect 185 72 191 74
rect 112 68 118 70
rect 185 70 187 72
rect 189 70 191 72
rect 185 68 191 70
<< nmos >>
rect -26 22 -24 31
rect -16 25 -14 31
rect -6 25 -4 31
rect 14 20 16 29
rect 27 18 29 29
rect 34 18 36 29
rect 54 22 56 31
rect 70 17 72 26
rect 80 17 82 26
rect 90 14 92 26
rect 97 14 99 26
rect 118 20 120 29
rect 131 18 133 29
rect 138 18 140 29
rect 158 22 160 31
rect 174 17 176 26
rect 184 17 186 26
rect 194 14 196 26
rect 201 14 203 26
<< pmos >>
rect -26 43 -24 61
rect -13 50 -11 71
rect -6 50 -4 71
rect 14 44 16 62
rect 24 51 26 64
rect 34 51 36 64
rect 62 44 64 71
rect 78 44 80 62
rect 88 44 90 62
rect 98 44 100 71
rect 118 44 120 62
rect 128 51 130 64
rect 138 51 140 64
rect 166 44 168 71
rect 182 44 184 62
rect 192 44 194 62
rect 202 44 204 71
<< polyct0 >>
rect -24 36 -22 38
rect 16 36 18 38
rect 86 36 88 38
rect 96 37 98 39
rect 120 36 122 38
rect 190 36 192 38
rect 200 37 202 39
<< polyct1 >>
rect -4 43 -2 45
rect -14 36 -12 38
rect 36 44 38 46
rect 49 44 51 46
rect 26 36 28 38
rect 140 44 142 46
rect 153 44 155 46
rect 65 31 67 33
rect 130 36 132 38
rect 169 31 171 33
<< ndifct0 >>
rect -11 27 -9 29
rect -20 14 -18 16
rect 49 27 51 29
rect 39 20 41 22
rect 63 19 65 21
rect -1 14 1 16
rect 75 22 77 24
rect 153 27 155 29
rect 143 20 145 22
rect 167 19 169 21
rect 179 22 181 24
<< ndifct1 >>
rect -31 27 -29 29
rect 9 22 11 24
rect 85 20 87 22
rect 20 10 22 12
rect 113 22 115 24
rect 103 10 105 12
rect 189 20 191 22
rect 124 10 126 12
rect 207 10 209 12
<< ntiect1 >>
rect -30 70 -28 72
rect 10 70 12 72
rect 83 70 85 72
rect 114 70 116 72
rect 187 70 189 72
<< ptiect1 >>
rect -30 10 -28 12
rect 10 10 12 12
rect 50 10 52 12
rect 114 10 116 12
rect 154 10 156 12
<< pdifct0 >>
rect -20 67 -18 69
rect -1 60 1 62
rect 19 58 21 60
rect 29 60 31 62
rect 29 53 31 55
rect 39 60 41 62
rect 57 46 59 48
rect 67 67 69 69
rect 67 60 69 62
rect 83 53 85 55
rect 83 46 85 48
rect 103 61 105 63
rect 123 58 125 60
rect 133 60 135 62
rect 133 53 135 55
rect 143 60 145 62
rect 161 46 163 48
rect 171 67 173 69
rect 171 60 173 62
rect 187 53 189 55
rect 187 46 189 48
rect 207 61 209 63
<< pdifct1 >>
rect -31 57 -29 59
rect -31 50 -29 52
rect 9 53 11 55
rect 9 46 11 48
rect 93 53 95 55
rect 113 53 115 55
rect 113 46 115 48
rect 197 53 199 55
<< alu0 >>
rect -22 67 -20 69
rect -18 67 -16 69
rect -22 66 -16 67
rect -14 62 3 63
rect -14 60 -1 62
rect 1 60 3 62
rect -14 59 3 60
rect 17 60 23 69
rect -29 48 -28 59
rect -14 55 -10 59
rect 17 58 19 60
rect 21 58 23 60
rect 17 57 23 58
rect 28 62 32 64
rect 28 60 29 62
rect 31 60 32 62
rect -25 51 -10 55
rect -25 38 -21 51
rect 28 55 32 60
rect 37 62 43 69
rect 66 67 67 69
rect 69 67 70 69
rect 37 60 39 62
rect 41 60 43 62
rect 37 59 43 60
rect 66 62 70 67
rect 66 60 67 62
rect 69 60 70 62
rect 66 58 70 60
rect 74 63 107 64
rect 74 61 103 63
rect 105 61 107 63
rect 74 60 107 61
rect 121 60 127 69
rect 28 54 29 55
rect 15 53 29 54
rect 31 53 32 55
rect 15 50 32 53
rect -6 42 0 43
rect -25 36 -24 38
rect -22 36 -21 38
rect -25 30 -21 36
rect -25 29 -7 30
rect -25 27 -11 29
rect -9 27 -7 29
rect -25 26 -7 27
rect 15 38 19 50
rect 74 49 78 60
rect 121 58 123 60
rect 125 58 127 60
rect 121 57 127 58
rect 132 62 136 64
rect 132 60 133 62
rect 135 60 136 62
rect 55 48 78 49
rect 55 46 57 48
rect 59 46 78 48
rect 55 45 78 46
rect 55 39 59 45
rect 15 36 16 38
rect 18 36 19 38
rect 15 31 19 36
rect 15 27 27 31
rect 11 24 12 26
rect 23 23 27 27
rect 48 35 59 39
rect 48 29 52 35
rect 74 39 78 45
rect 82 55 86 57
rect 82 53 83 55
rect 85 53 86 55
rect 82 48 86 53
rect 82 46 83 48
rect 85 47 86 48
rect 85 46 98 47
rect 82 43 98 46
rect 94 41 98 43
rect 94 39 99 41
rect 74 38 90 39
rect 74 36 86 38
rect 88 36 90 38
rect 74 35 90 36
rect 94 37 96 39
rect 98 37 99 39
rect 94 35 99 37
rect 48 27 49 29
rect 51 27 52 29
rect 48 25 52 27
rect 94 31 98 35
rect 74 27 98 31
rect 74 24 78 27
rect 23 22 43 23
rect 74 22 75 24
rect 77 22 78 24
rect 23 20 39 22
rect 41 20 43 22
rect 23 19 43 20
rect 61 21 67 22
rect 61 19 63 21
rect 65 19 67 21
rect 74 20 78 22
rect 132 55 136 60
rect 141 62 147 69
rect 170 67 171 69
rect 173 67 174 69
rect 141 60 143 62
rect 145 60 147 62
rect 141 59 147 60
rect 170 62 174 67
rect 170 60 171 62
rect 173 60 174 62
rect 170 58 174 60
rect 178 63 211 64
rect 178 61 207 63
rect 209 61 211 63
rect 178 60 211 61
rect 132 54 133 55
rect 119 53 133 54
rect 135 53 136 55
rect 119 50 136 53
rect 119 38 123 50
rect 178 49 182 60
rect 159 48 182 49
rect 159 46 161 48
rect 163 46 182 48
rect 159 45 182 46
rect 159 39 163 45
rect 119 36 120 38
rect 122 36 123 38
rect 119 31 123 36
rect 119 27 131 31
rect 115 24 116 26
rect -22 16 -16 17
rect -22 14 -20 16
rect -18 14 -16 16
rect -22 13 -16 14
rect -3 16 3 17
rect -3 14 -1 16
rect 1 14 3 16
rect -3 13 3 14
rect 61 13 67 19
rect 127 23 131 27
rect 152 35 163 39
rect 152 29 156 35
rect 178 39 182 45
rect 186 55 190 57
rect 186 53 187 55
rect 189 53 190 55
rect 186 48 190 53
rect 186 46 187 48
rect 189 47 190 48
rect 189 46 202 47
rect 186 43 202 46
rect 198 41 202 43
rect 198 39 203 41
rect 178 38 194 39
rect 178 36 190 38
rect 192 36 194 38
rect 178 35 194 36
rect 198 37 200 39
rect 202 37 203 39
rect 198 35 203 37
rect 152 27 153 29
rect 155 27 156 29
rect 152 25 156 27
rect 198 31 202 35
rect 178 27 202 31
rect 178 24 182 27
rect 127 22 147 23
rect 178 22 179 24
rect 181 22 182 24
rect 127 20 143 22
rect 145 20 147 22
rect 127 19 147 20
rect 165 21 171 22
rect 165 19 167 21
rect 169 19 171 21
rect 178 20 182 22
rect 165 13 171 19
<< via1 >>
rect 0 49 2 51
rect 8 49 10 51
rect 40 51 42 53
rect 0 36 2 38
rect 49 51 51 53
rect 32 27 34 29
rect 104 44 106 46
rect 57 27 59 29
rect 144 51 146 53
rect 112 36 114 38
rect 135 44 137 46
rect 153 51 155 53
rect 136 27 138 29
rect 161 27 163 29
<< labels >>
rlabel alu0 50 32 50 32 6 bn
rlabel alu0 96 37 96 37 6 an
rlabel alu1 65 33 65 33 6 a
rlabel alu1 77 9 77 9 6 vss
rlabel alu1 77 73 77 73 6 vdd
rlabel alu1 41 53 41 53 6 b
rlabel alu1 25 73 25 73 6 vdd
rlabel alu1 25 37 25 37 6 a
rlabel alu1 25 9 25 9 6 vss
rlabel alu0 17 40 17 40 6 zn
rlabel alu1 129 9 129 9 6 vss
rlabel alu1 129 73 129 73 6 vdd
rlabel alu1 209 33 209 33 1 sum
rlabel alu1 181 73 181 73 6 vdd
rlabel alu1 181 9 181 9 6 vss
rlabel alu1 105 33 105 33 1 s
rlabel alu1 129 36 129 36 1 cin
rlabel alu1 17 21 17 21 1 co
rlabel alu0 121 39 121 39 1 zn_1
rlabel alu0 154 32 154 32 1 bn_1
rlabel alu0 180 24 180 24 1 an_1
rlabel alu1 -15 73 -15 73 6 vdd
rlabel alu1 -15 9 -15 9 6 vss
rlabel alu1 121 21 121 21 1 c1
rlabel alu1 -31 41 -31 41 1 cout
rlabel alu0 -6 61 -6 61 1 zn_2
<< end >>
