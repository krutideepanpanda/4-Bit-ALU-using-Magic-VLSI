magic
tech scmos
timestamp 1636300124
<< ab >>
rect 44 446 50 451
rect 148 446 154 451
rect -31 445 217 446
rect -31 444 131 445
rect -31 441 -14 444
rect -10 441 27 444
rect -31 440 27 441
rect 31 443 131 444
rect 31 440 80 443
rect 82 441 131 443
rect 135 443 217 445
rect 135 441 183 443
rect 82 440 183 441
rect 187 440 217 443
rect -31 414 217 440
rect -31 382 49 414
rect 50 382 153 414
rect 154 382 217 414
rect -31 380 217 382
rect -31 376 -14 380
rect -9 376 26 380
rect 30 376 79 380
rect 83 376 130 380
rect 134 376 183 380
rect 187 376 217 380
rect -31 372 217 376
rect -31 368 -14 372
rect -9 368 26 372
rect 30 368 79 372
rect 83 368 130 372
rect 134 368 183 372
rect 187 368 217 372
rect -31 366 217 368
rect -31 334 49 366
rect 50 334 153 366
rect 154 334 217 366
rect -31 308 217 334
rect -31 307 27 308
rect -31 304 -14 307
rect -10 304 27 307
rect 31 305 80 308
rect 82 307 183 308
rect 82 305 131 307
rect 31 304 131 305
rect -31 303 131 304
rect 135 305 183 307
rect 187 305 217 308
rect 135 303 217 305
rect -31 301 217 303
rect -31 300 131 301
rect -31 297 -14 300
rect -10 297 27 300
rect -31 296 27 297
rect 31 299 131 300
rect 31 296 80 299
rect 82 297 131 299
rect 135 299 217 301
rect 135 297 183 299
rect 82 296 183 297
rect 187 296 217 299
rect -31 270 217 296
rect -31 238 49 270
rect 50 238 153 270
rect 154 238 217 270
rect -31 236 217 238
rect -31 232 -14 236
rect -9 232 26 236
rect 30 232 79 236
rect 83 232 130 236
rect 134 232 183 236
rect 187 232 217 236
rect -31 228 217 232
rect -31 224 -14 228
rect -9 224 26 228
rect 30 224 79 228
rect 83 224 130 228
rect 134 224 183 228
rect 187 224 217 228
rect -31 222 217 224
rect -31 190 49 222
rect 50 190 153 222
rect 154 190 217 222
rect -31 164 217 190
rect -31 163 27 164
rect -31 160 -14 163
rect -10 160 27 163
rect 31 161 80 164
rect 82 163 183 164
rect 82 161 131 163
rect 31 160 131 161
rect -31 159 131 160
rect 135 161 183 163
rect 187 161 217 164
rect 135 159 217 161
rect -31 158 217 159
rect 226 444 266 446
rect 226 440 244 444
rect 248 440 266 444
rect 226 431 266 440
rect 226 429 237 431
rect 239 429 253 431
rect 255 429 266 431
rect 226 415 266 429
rect 226 413 261 415
rect 263 413 266 415
rect 226 412 266 413
rect 226 410 253 412
rect 255 410 266 412
rect 226 395 266 410
rect 226 393 240 395
rect 242 393 266 395
rect 226 380 266 393
rect 226 376 244 380
rect 248 376 266 380
rect 226 372 266 376
rect 226 368 244 372
rect 248 368 266 372
rect 226 355 266 368
rect 226 353 240 355
rect 242 353 266 355
rect 226 338 266 353
rect 226 336 253 338
rect 255 336 266 338
rect 226 335 266 336
rect 226 333 261 335
rect 263 333 266 335
rect 226 319 266 333
rect 226 317 237 319
rect 239 317 253 319
rect 255 317 266 319
rect 226 308 266 317
rect 226 304 244 308
rect 248 304 266 308
rect 226 300 266 304
rect 226 296 244 300
rect 248 296 266 300
rect 226 287 266 296
rect 226 285 237 287
rect 239 285 253 287
rect 255 285 266 287
rect 226 271 266 285
rect 226 269 261 271
rect 263 269 266 271
rect 226 268 266 269
rect 226 266 253 268
rect 255 266 266 268
rect 226 251 266 266
rect 226 249 240 251
rect 242 249 266 251
rect 226 236 266 249
rect 226 232 244 236
rect 248 232 266 236
rect 226 228 266 232
rect 226 224 244 228
rect 248 224 266 228
rect 226 211 266 224
rect 226 209 240 211
rect 242 209 266 211
rect 226 194 266 209
rect 226 192 253 194
rect 255 192 266 194
rect 226 191 266 192
rect 226 189 261 191
rect 263 189 266 191
rect 226 175 266 189
rect 226 173 237 175
rect 239 173 253 175
rect 255 173 266 175
rect 226 164 266 173
rect 226 160 244 164
rect 248 160 266 164
rect 226 158 266 160
rect 274 444 314 446
rect 274 441 292 444
rect 296 441 314 444
rect 274 424 314 441
rect 274 422 294 424
rect 296 422 314 424
rect 274 412 314 422
rect 274 410 301 412
rect 303 410 314 412
rect 274 407 314 410
rect 274 405 309 407
rect 311 405 314 407
rect 274 391 314 405
rect 274 389 284 391
rect 286 389 301 391
rect 303 389 314 391
rect 274 380 314 389
rect 274 376 292 380
rect 296 376 314 380
rect 274 372 314 376
rect 274 368 292 372
rect 296 368 314 372
rect 274 359 314 368
rect 274 357 284 359
rect 286 357 301 359
rect 303 357 314 359
rect 274 343 314 357
rect 274 341 309 343
rect 311 341 314 343
rect 274 338 314 341
rect 274 336 301 338
rect 303 336 314 338
rect 274 326 314 336
rect 274 324 294 326
rect 296 324 314 326
rect 274 307 314 324
rect 274 304 292 307
rect 296 304 314 307
rect 274 300 314 304
rect 274 297 292 300
rect 296 297 314 300
rect 274 280 314 297
rect 274 278 294 280
rect 296 278 314 280
rect 274 268 314 278
rect 274 266 301 268
rect 303 266 314 268
rect 274 263 314 266
rect 274 261 309 263
rect 311 261 314 263
rect 274 247 314 261
rect 274 245 284 247
rect 286 245 301 247
rect 303 245 314 247
rect 274 236 314 245
rect 274 232 292 236
rect 296 232 314 236
rect 274 228 314 232
rect 274 224 292 228
rect 296 224 314 228
rect 274 215 314 224
rect 274 213 284 215
rect 286 213 301 215
rect 303 213 314 215
rect 274 199 314 213
rect 274 197 309 199
rect 311 197 314 199
rect 274 194 314 197
rect 274 192 301 194
rect 303 192 314 194
rect 274 182 314 192
rect 274 180 294 182
rect 296 180 314 182
rect 274 163 314 180
rect 274 160 292 163
rect 296 160 314 163
rect 274 158 314 160
rect 323 443 387 446
rect 323 441 354 443
rect 356 441 387 443
rect 323 433 387 441
rect 323 429 349 433
rect 351 429 387 433
rect 323 423 387 429
rect 323 421 374 423
rect 376 421 387 423
rect 323 419 354 421
rect 356 419 387 421
rect 323 418 387 419
rect 323 416 382 418
rect 384 416 387 418
rect 323 415 387 416
rect 323 413 326 415
rect 328 413 366 415
rect 370 413 387 415
rect 323 411 358 413
rect 360 411 387 413
rect 323 409 334 411
rect 336 409 342 411
rect 344 409 387 411
rect 323 407 387 409
rect 323 405 350 407
rect 352 406 387 407
rect 352 405 370 406
rect 323 404 370 405
rect 372 404 387 406
rect 323 399 387 404
rect 323 397 374 399
rect 376 397 387 399
rect 323 395 387 397
rect 323 392 349 395
rect 353 392 387 395
rect 323 391 387 392
rect 323 389 334 391
rect 336 389 382 391
rect 384 389 387 391
rect 323 379 387 389
rect 323 377 354 379
rect 356 377 387 379
rect 323 371 387 377
rect 323 369 354 371
rect 356 369 387 371
rect 323 359 387 369
rect 323 357 334 359
rect 336 357 382 359
rect 384 357 387 359
rect 323 356 387 357
rect 323 353 349 356
rect 353 353 387 356
rect 323 351 387 353
rect 323 349 374 351
rect 376 349 387 351
rect 323 344 387 349
rect 323 343 370 344
rect 323 341 350 343
rect 352 342 370 343
rect 372 342 387 344
rect 352 341 387 342
rect 323 339 387 341
rect 323 337 334 339
rect 336 337 342 339
rect 344 337 387 339
rect 323 335 358 337
rect 360 335 387 337
rect 323 333 326 335
rect 328 333 366 335
rect 370 333 387 335
rect 323 332 387 333
rect 323 330 382 332
rect 384 330 387 332
rect 323 329 387 330
rect 323 327 354 329
rect 356 327 387 329
rect 323 325 374 327
rect 376 325 387 327
rect 323 319 387 325
rect 323 315 349 319
rect 351 315 387 319
rect 323 307 387 315
rect 323 305 354 307
rect 356 305 387 307
rect 323 299 387 305
rect 323 297 354 299
rect 356 297 387 299
rect 323 289 387 297
rect 323 285 349 289
rect 351 285 387 289
rect 323 279 387 285
rect 323 277 374 279
rect 376 277 387 279
rect 323 275 354 277
rect 356 275 387 277
rect 323 274 387 275
rect 323 272 382 274
rect 384 272 387 274
rect 323 271 387 272
rect 323 269 326 271
rect 328 269 366 271
rect 370 269 387 271
rect 323 267 358 269
rect 360 267 387 269
rect 323 265 334 267
rect 336 265 342 267
rect 344 265 387 267
rect 323 263 387 265
rect 323 261 350 263
rect 352 262 387 263
rect 352 261 370 262
rect 323 260 370 261
rect 372 260 387 262
rect 323 255 387 260
rect 323 253 374 255
rect 376 253 387 255
rect 323 251 387 253
rect 323 248 349 251
rect 353 248 387 251
rect 323 247 387 248
rect 323 245 334 247
rect 336 245 382 247
rect 384 245 387 247
rect 323 235 387 245
rect 323 233 354 235
rect 356 233 387 235
rect 323 227 387 233
rect 323 225 354 227
rect 356 225 387 227
rect 323 215 387 225
rect 323 213 334 215
rect 336 213 382 215
rect 384 213 387 215
rect 323 212 387 213
rect 323 209 349 212
rect 353 209 387 212
rect 323 207 387 209
rect 323 205 374 207
rect 376 205 387 207
rect 323 200 387 205
rect 323 199 370 200
rect 323 197 350 199
rect 352 198 370 199
rect 372 198 387 200
rect 352 197 387 198
rect 323 195 387 197
rect 323 193 334 195
rect 336 193 342 195
rect 344 193 387 195
rect 323 191 358 193
rect 360 191 387 193
rect 323 189 326 191
rect 328 189 366 191
rect 370 189 387 191
rect 323 188 387 189
rect 323 186 382 188
rect 384 186 387 188
rect 323 185 387 186
rect 323 183 354 185
rect 356 183 387 185
rect 323 181 374 183
rect 376 181 387 183
rect 323 175 387 181
rect 323 171 349 175
rect 351 171 387 175
rect 323 163 387 171
rect 323 161 354 163
rect 356 161 387 163
rect 323 158 387 161
rect 397 443 461 446
rect 397 441 428 443
rect 430 441 461 443
rect 397 433 461 441
rect 397 429 423 433
rect 425 429 461 433
rect 397 423 461 429
rect 397 421 448 423
rect 450 421 461 423
rect 397 419 428 421
rect 430 419 461 421
rect 397 418 461 419
rect 397 416 456 418
rect 458 416 461 418
rect 397 415 461 416
rect 397 413 400 415
rect 402 413 440 415
rect 442 413 461 415
rect 397 411 432 413
rect 434 411 461 413
rect 397 409 408 411
rect 410 409 416 411
rect 418 409 461 411
rect 397 407 461 409
rect 397 405 424 407
rect 426 406 461 407
rect 426 405 444 406
rect 397 404 444 405
rect 446 404 461 406
rect 397 399 461 404
rect 397 397 448 399
rect 450 397 461 399
rect 397 395 461 397
rect 397 392 423 395
rect 427 392 461 395
rect 397 391 461 392
rect 397 389 408 391
rect 410 389 456 391
rect 458 389 461 391
rect 397 379 461 389
rect 397 377 428 379
rect 430 377 461 379
rect 397 371 461 377
rect 397 369 428 371
rect 430 369 461 371
rect 397 359 461 369
rect 397 357 408 359
rect 410 357 456 359
rect 458 357 461 359
rect 397 356 461 357
rect 397 353 423 356
rect 427 353 461 356
rect 397 351 461 353
rect 397 349 448 351
rect 450 349 461 351
rect 397 344 461 349
rect 397 343 444 344
rect 397 341 424 343
rect 426 342 444 343
rect 446 342 461 344
rect 426 341 461 342
rect 397 339 461 341
rect 397 337 408 339
rect 410 337 416 339
rect 418 337 461 339
rect 397 335 432 337
rect 434 335 461 337
rect 397 333 400 335
rect 402 333 440 335
rect 442 333 461 335
rect 397 332 461 333
rect 397 330 456 332
rect 458 330 461 332
rect 397 329 461 330
rect 397 327 428 329
rect 430 327 461 329
rect 397 325 448 327
rect 450 325 461 327
rect 397 319 461 325
rect 397 315 423 319
rect 425 315 461 319
rect 397 307 461 315
rect 397 305 428 307
rect 430 305 461 307
rect 397 299 461 305
rect 397 297 428 299
rect 430 297 461 299
rect 397 289 461 297
rect 397 285 423 289
rect 425 285 461 289
rect 397 279 461 285
rect 397 277 448 279
rect 450 277 461 279
rect 397 275 428 277
rect 430 275 461 277
rect 397 274 461 275
rect 397 272 456 274
rect 458 272 461 274
rect 397 271 461 272
rect 397 269 400 271
rect 402 269 440 271
rect 442 269 461 271
rect 397 267 432 269
rect 434 267 461 269
rect 397 265 408 267
rect 410 265 416 267
rect 418 265 461 267
rect 397 263 461 265
rect 397 261 424 263
rect 426 262 461 263
rect 426 261 444 262
rect 397 260 444 261
rect 446 260 461 262
rect 397 255 461 260
rect 397 253 448 255
rect 450 253 461 255
rect 397 251 461 253
rect 397 248 423 251
rect 427 248 461 251
rect 397 247 461 248
rect 397 245 408 247
rect 410 245 456 247
rect 458 245 461 247
rect 397 235 461 245
rect 397 233 428 235
rect 430 233 461 235
rect 397 227 461 233
rect 397 225 428 227
rect 430 225 461 227
rect 397 215 461 225
rect 397 213 408 215
rect 410 213 456 215
rect 458 213 461 215
rect 397 212 461 213
rect 397 209 423 212
rect 427 209 461 212
rect 397 207 461 209
rect 397 205 448 207
rect 450 205 461 207
rect 397 200 461 205
rect 397 199 444 200
rect 397 197 424 199
rect 426 198 444 199
rect 446 198 461 200
rect 426 197 461 198
rect 397 195 461 197
rect 397 193 408 195
rect 410 193 416 195
rect 418 193 461 195
rect 397 191 432 193
rect 434 191 461 193
rect 397 189 400 191
rect 402 189 440 191
rect 442 189 461 191
rect 397 188 461 189
rect 397 186 456 188
rect 458 186 461 188
rect 397 185 461 186
rect 397 183 428 185
rect 430 183 461 185
rect 397 181 448 183
rect 450 181 461 183
rect 397 175 461 181
rect 397 171 423 175
rect 425 171 461 175
rect 397 163 461 171
rect 397 161 428 163
rect 430 161 461 163
rect 397 158 461 161
rect 471 443 535 446
rect 471 441 502 443
rect 504 441 535 443
rect 471 433 535 441
rect 471 429 497 433
rect 499 429 535 433
rect 471 423 535 429
rect 471 421 522 423
rect 524 421 535 423
rect 471 419 502 421
rect 504 419 535 421
rect 471 418 535 419
rect 471 416 530 418
rect 532 416 535 418
rect 471 415 535 416
rect 471 413 474 415
rect 476 413 514 415
rect 516 413 535 415
rect 471 412 506 413
rect 471 410 474 412
rect 476 411 506 412
rect 508 411 535 413
rect 476 410 482 411
rect 471 409 482 410
rect 484 409 490 411
rect 492 409 535 411
rect 471 407 535 409
rect 471 405 498 407
rect 500 406 535 407
rect 500 405 518 406
rect 471 404 518 405
rect 520 404 535 406
rect 471 399 535 404
rect 471 397 522 399
rect 524 397 535 399
rect 471 395 535 397
rect 471 392 497 395
rect 501 392 535 395
rect 471 391 535 392
rect 471 389 482 391
rect 484 389 530 391
rect 532 389 535 391
rect 471 379 535 389
rect 471 377 502 379
rect 504 377 535 379
rect 471 371 535 377
rect 471 369 502 371
rect 504 369 535 371
rect 471 359 535 369
rect 471 357 482 359
rect 484 357 530 359
rect 532 357 535 359
rect 471 356 535 357
rect 471 353 497 356
rect 501 353 535 356
rect 471 351 535 353
rect 471 349 522 351
rect 524 349 535 351
rect 471 344 535 349
rect 471 343 518 344
rect 471 341 498 343
rect 500 342 518 343
rect 520 342 535 344
rect 500 341 535 342
rect 471 339 535 341
rect 471 338 482 339
rect 471 336 474 338
rect 476 337 482 338
rect 484 337 490 339
rect 492 337 535 339
rect 476 336 506 337
rect 471 335 506 336
rect 508 335 535 337
rect 471 333 474 335
rect 476 333 514 335
rect 516 333 535 335
rect 471 332 535 333
rect 471 330 530 332
rect 532 330 535 332
rect 471 329 535 330
rect 471 327 502 329
rect 504 327 535 329
rect 471 325 522 327
rect 524 325 535 327
rect 471 319 535 325
rect 471 315 497 319
rect 499 315 535 319
rect 471 307 535 315
rect 471 305 502 307
rect 504 305 535 307
rect 471 299 535 305
rect 471 297 502 299
rect 504 297 535 299
rect 471 289 535 297
rect 471 285 497 289
rect 499 285 535 289
rect 471 279 535 285
rect 471 277 522 279
rect 524 277 535 279
rect 471 275 502 277
rect 504 275 535 277
rect 471 274 535 275
rect 471 272 530 274
rect 532 272 535 274
rect 471 271 535 272
rect 471 269 474 271
rect 476 269 514 271
rect 516 269 535 271
rect 471 268 506 269
rect 471 266 474 268
rect 476 267 506 268
rect 508 267 535 269
rect 476 266 482 267
rect 471 265 482 266
rect 484 265 490 267
rect 492 265 535 267
rect 471 263 535 265
rect 471 261 498 263
rect 500 262 535 263
rect 500 261 518 262
rect 471 260 518 261
rect 520 260 535 262
rect 471 255 535 260
rect 471 253 522 255
rect 524 253 535 255
rect 471 251 535 253
rect 471 248 497 251
rect 501 248 535 251
rect 471 247 535 248
rect 471 245 482 247
rect 484 245 530 247
rect 532 245 535 247
rect 471 235 535 245
rect 471 233 502 235
rect 504 233 535 235
rect 471 227 535 233
rect 471 225 502 227
rect 504 225 535 227
rect 471 215 535 225
rect 471 213 482 215
rect 484 213 530 215
rect 532 213 535 215
rect 471 212 535 213
rect 471 209 497 212
rect 501 209 535 212
rect 471 207 535 209
rect 471 205 522 207
rect 524 205 535 207
rect 471 200 535 205
rect 471 199 518 200
rect 471 197 498 199
rect 500 198 518 199
rect 520 198 535 200
rect 500 197 535 198
rect 471 195 535 197
rect 471 194 482 195
rect 471 192 474 194
rect 476 193 482 194
rect 484 193 490 195
rect 492 193 535 195
rect 476 192 506 193
rect 471 191 506 192
rect 508 191 535 193
rect 471 189 474 191
rect 476 189 514 191
rect 516 189 535 191
rect 471 188 535 189
rect 471 186 530 188
rect 532 186 535 188
rect 471 185 535 186
rect 471 183 502 185
rect 504 183 535 185
rect 471 181 522 183
rect 524 181 535 183
rect 471 175 535 181
rect 471 171 497 175
rect 499 171 535 175
rect 471 163 535 171
rect 471 161 502 163
rect 504 161 535 163
rect 471 158 535 161
<< nwell >>
rect -37 334 540 414
rect -37 190 540 270
<< pwell >>
rect -37 414 540 451
rect -37 270 540 334
rect -37 158 540 190
<< poly >>
rect -22 429 -20 434
rect -12 426 -10 431
rect -2 426 0 431
rect 18 431 20 435
rect 31 433 33 438
rect 38 433 40 438
rect 61 442 86 444
rect 61 434 63 442
rect 74 434 76 438
rect 84 434 86 442
rect 94 437 96 442
rect 101 437 103 442
rect 58 432 63 434
rect 58 429 60 432
rect -22 417 -20 420
rect -12 417 -10 420
rect -22 415 -16 417
rect -22 413 -20 415
rect -18 413 -16 415
rect -22 411 -16 413
rect -12 415 -6 417
rect -12 413 -10 415
rect -8 413 -6 415
rect -12 411 -6 413
rect -22 408 -20 411
rect -9 401 -7 411
rect -2 410 0 420
rect 18 417 20 422
rect 31 417 33 422
rect 18 415 24 417
rect 18 413 20 415
rect 22 413 24 415
rect 18 411 24 413
rect 28 415 34 417
rect 28 413 30 415
rect 32 413 34 415
rect 28 411 34 413
rect -2 408 4 410
rect -2 406 0 408
rect 2 406 4 408
rect 18 407 20 411
rect -2 404 4 406
rect -2 401 0 404
rect -22 385 -20 390
rect 28 400 30 411
rect 38 409 40 422
rect 122 431 124 435
rect 135 433 137 438
rect 142 433 144 438
rect 165 442 190 444
rect 165 434 167 442
rect 178 434 180 438
rect 188 434 190 442
rect 198 437 200 442
rect 205 437 207 442
rect 74 422 76 425
rect 67 420 76 422
rect 84 421 86 425
rect 94 422 96 425
rect 58 412 60 420
rect 67 418 69 420
rect 71 418 76 420
rect 67 416 76 418
rect 92 420 96 422
rect 92 417 94 420
rect 74 412 76 416
rect 88 415 94 417
rect 101 416 103 425
rect 162 432 167 434
rect 162 429 164 432
rect 122 417 124 422
rect 135 417 137 422
rect 88 413 90 415
rect 92 413 94 415
rect 55 410 68 412
rect 74 410 84 412
rect 88 411 94 413
rect 55 409 57 410
rect 38 407 44 409
rect 38 405 40 407
rect 42 405 44 407
rect 38 403 44 405
rect 51 407 57 409
rect 66 407 68 410
rect 82 407 84 410
rect 92 407 94 411
rect 98 414 104 416
rect 98 412 100 414
rect 102 412 104 414
rect 98 410 104 412
rect 102 407 104 410
rect 122 415 128 417
rect 122 413 124 415
rect 126 413 128 415
rect 122 411 128 413
rect 132 415 138 417
rect 132 413 134 415
rect 136 413 138 415
rect 132 411 138 413
rect 122 407 124 411
rect 51 405 53 407
rect 55 405 57 407
rect 51 403 57 405
rect 38 400 40 403
rect 18 385 20 389
rect 28 382 30 387
rect 38 382 40 387
rect -9 376 -7 380
rect -2 376 0 380
rect 82 385 84 389
rect 92 385 94 389
rect 66 376 68 380
rect 132 400 134 411
rect 142 409 144 422
rect 235 433 237 438
rect 242 433 244 438
rect 359 442 378 444
rect 178 422 180 425
rect 171 420 180 422
rect 188 421 190 425
rect 198 422 200 425
rect 162 412 164 420
rect 171 418 173 420
rect 175 418 180 420
rect 171 416 180 418
rect 196 420 200 422
rect 196 417 198 420
rect 178 412 180 416
rect 192 415 198 417
rect 205 416 207 425
rect 255 431 257 435
rect 332 434 334 439
rect 342 434 344 439
rect 349 434 351 439
rect 359 434 361 442
rect 366 434 368 438
rect 283 426 285 431
rect 293 426 295 431
rect 303 429 305 434
rect 192 413 194 415
rect 196 413 198 415
rect 159 410 172 412
rect 178 410 188 412
rect 192 411 198 413
rect 159 409 161 410
rect 142 407 148 409
rect 142 405 144 407
rect 146 405 148 407
rect 142 403 148 405
rect 155 407 161 409
rect 170 407 172 410
rect 186 407 188 410
rect 196 407 198 411
rect 202 414 208 416
rect 202 412 204 414
rect 206 412 208 414
rect 202 410 208 412
rect 206 407 208 410
rect 235 409 237 422
rect 242 417 244 422
rect 255 417 257 422
rect 376 432 378 442
rect 433 442 452 444
rect 406 434 408 439
rect 416 434 418 439
rect 423 434 425 439
rect 433 434 435 442
rect 440 434 442 438
rect 332 422 334 425
rect 331 420 337 422
rect 241 415 247 417
rect 241 413 243 415
rect 245 413 247 415
rect 241 411 247 413
rect 251 415 257 417
rect 251 413 253 415
rect 255 413 257 415
rect 251 411 257 413
rect 231 407 237 409
rect 155 405 157 407
rect 159 405 161 407
rect 155 403 161 405
rect 142 400 144 403
rect 122 385 124 389
rect 132 382 134 387
rect 142 382 144 387
rect 102 376 104 380
rect 186 385 188 389
rect 196 385 198 389
rect 170 376 172 380
rect 231 405 233 407
rect 235 405 237 407
rect 231 403 237 405
rect 235 400 237 403
rect 245 400 247 411
rect 255 407 257 411
rect 283 410 285 420
rect 293 417 295 420
rect 303 417 305 420
rect 289 415 295 417
rect 289 413 291 415
rect 293 413 295 415
rect 289 411 295 413
rect 299 415 305 417
rect 331 418 333 420
rect 335 418 337 420
rect 331 416 337 418
rect 299 413 301 415
rect 303 413 305 415
rect 299 411 305 413
rect 279 408 285 410
rect 279 406 281 408
rect 283 406 285 408
rect 279 404 285 406
rect 283 401 285 404
rect 290 401 292 411
rect 303 408 305 411
rect 235 382 237 387
rect 245 382 247 387
rect 255 385 257 389
rect 206 376 208 380
rect 332 398 334 416
rect 342 412 344 426
rect 349 423 351 426
rect 349 421 355 423
rect 349 419 351 421
rect 353 419 355 421
rect 349 417 355 419
rect 359 413 361 426
rect 339 410 345 412
rect 339 408 341 410
rect 343 408 345 410
rect 339 406 345 408
rect 349 411 361 413
rect 366 422 368 426
rect 366 420 372 422
rect 366 418 368 420
rect 370 418 372 420
rect 366 411 372 418
rect 303 385 305 390
rect 283 376 285 380
rect 290 376 292 380
rect 342 396 344 406
rect 349 396 351 411
rect 356 405 362 407
rect 356 403 358 405
rect 360 403 362 405
rect 356 401 362 403
rect 359 396 361 401
rect 366 396 368 411
rect 376 408 378 426
rect 450 432 452 442
rect 507 442 526 444
rect 480 434 482 439
rect 490 434 492 439
rect 497 434 499 439
rect 507 434 509 442
rect 514 434 516 438
rect 406 422 408 425
rect 405 420 411 422
rect 405 418 407 420
rect 409 418 411 420
rect 405 416 411 418
rect 376 397 378 400
rect 406 398 408 416
rect 416 412 418 426
rect 423 423 425 426
rect 423 421 429 423
rect 423 419 425 421
rect 427 419 429 421
rect 423 417 429 419
rect 433 413 435 426
rect 413 410 419 412
rect 413 408 415 410
rect 417 408 419 410
rect 413 406 419 408
rect 423 411 435 413
rect 440 417 442 426
rect 440 415 446 417
rect 440 413 442 415
rect 444 413 446 415
rect 440 411 446 413
rect 376 395 385 397
rect 379 393 381 395
rect 383 393 385 395
rect 379 391 385 393
rect 416 396 418 406
rect 423 396 425 411
rect 430 405 436 407
rect 430 403 432 405
rect 434 403 436 405
rect 430 401 436 403
rect 433 396 435 401
rect 440 396 442 411
rect 450 408 452 426
rect 524 432 526 442
rect 480 422 482 425
rect 479 420 485 422
rect 479 418 481 420
rect 483 418 485 420
rect 479 416 485 418
rect 450 397 452 400
rect 480 398 482 416
rect 490 412 492 426
rect 497 423 499 426
rect 497 421 503 423
rect 497 419 499 421
rect 501 419 503 421
rect 497 417 503 419
rect 507 413 509 426
rect 487 410 493 412
rect 487 408 489 410
rect 491 408 493 410
rect 487 406 493 408
rect 497 411 509 413
rect 514 417 516 426
rect 514 415 520 417
rect 514 413 516 415
rect 518 413 520 415
rect 514 411 520 413
rect 450 395 459 397
rect 453 393 455 395
rect 457 393 459 395
rect 453 391 459 393
rect 490 396 492 406
rect 497 396 499 411
rect 504 405 510 407
rect 504 403 506 405
rect 508 403 510 405
rect 504 401 510 403
rect 507 396 509 401
rect 514 396 516 411
rect 524 408 526 426
rect 524 397 526 400
rect 524 395 533 397
rect 527 393 529 395
rect 531 393 533 395
rect 527 391 533 393
rect 332 376 334 380
rect 342 376 344 380
rect 349 376 351 380
rect 359 376 361 380
rect 366 376 368 380
rect 406 376 408 380
rect 416 376 418 380
rect 423 376 425 380
rect 433 376 435 380
rect 440 376 442 380
rect 480 376 482 380
rect 490 376 492 380
rect 497 376 499 380
rect 507 376 509 380
rect 514 376 516 380
rect -9 368 -7 372
rect -2 368 0 372
rect -22 358 -20 363
rect 66 368 68 372
rect 18 359 20 363
rect 28 361 30 366
rect 38 361 40 366
rect -22 337 -20 340
rect -9 337 -7 347
rect -2 344 0 347
rect -2 342 4 344
rect -2 340 0 342
rect 2 340 4 342
rect -2 338 4 340
rect -22 335 -16 337
rect -22 333 -20 335
rect -18 333 -16 335
rect -22 331 -16 333
rect -12 335 -6 337
rect -12 333 -10 335
rect -8 333 -6 335
rect -12 331 -6 333
rect -22 328 -20 331
rect -12 328 -10 331
rect -2 328 0 338
rect 18 337 20 341
rect 28 337 30 348
rect 38 345 40 348
rect 38 343 44 345
rect 38 341 40 343
rect 42 341 44 343
rect 38 339 44 341
rect 51 343 57 345
rect 51 341 53 343
rect 55 341 57 343
rect 102 368 104 372
rect 82 359 84 363
rect 92 359 94 363
rect 170 368 172 372
rect 122 359 124 363
rect 132 361 134 366
rect 142 361 144 366
rect 51 339 57 341
rect 18 335 24 337
rect 18 333 20 335
rect 22 333 24 335
rect 18 331 24 333
rect 28 335 34 337
rect 28 333 30 335
rect 32 333 34 335
rect 28 331 34 333
rect 18 326 20 331
rect 31 326 33 331
rect 38 326 40 339
rect 55 338 57 339
rect 66 338 68 341
rect 82 338 84 341
rect 55 336 68 338
rect 74 336 84 338
rect 92 337 94 341
rect 102 338 104 341
rect 58 328 60 336
rect 74 332 76 336
rect 67 330 76 332
rect 88 335 94 337
rect 88 333 90 335
rect 92 333 94 335
rect 88 331 94 333
rect 98 336 104 338
rect 98 334 100 336
rect 102 334 104 336
rect 98 332 104 334
rect 122 337 124 341
rect 132 337 134 348
rect 142 345 144 348
rect 142 343 148 345
rect 142 341 144 343
rect 146 341 148 343
rect 142 339 148 341
rect 155 343 161 345
rect 155 341 157 343
rect 159 341 161 343
rect 206 368 208 372
rect 186 359 188 363
rect 196 359 198 363
rect 283 368 285 372
rect 290 368 292 372
rect 235 361 237 366
rect 245 361 247 366
rect 255 359 257 363
rect 235 345 237 348
rect 231 343 237 345
rect 231 341 233 343
rect 235 341 237 343
rect 155 339 161 341
rect 122 335 128 337
rect 122 333 124 335
rect 126 333 128 335
rect 67 328 69 330
rect 71 328 76 330
rect -22 314 -20 319
rect -12 317 -10 322
rect -2 317 0 322
rect 18 313 20 317
rect 67 326 76 328
rect 92 328 94 331
rect 74 323 76 326
rect 84 323 86 327
rect 92 326 96 328
rect 94 323 96 326
rect 101 323 103 332
rect 122 331 128 333
rect 132 335 138 337
rect 132 333 134 335
rect 136 333 138 335
rect 132 331 138 333
rect 122 326 124 331
rect 135 326 137 331
rect 142 326 144 339
rect 159 338 161 339
rect 170 338 172 341
rect 186 338 188 341
rect 159 336 172 338
rect 178 336 188 338
rect 196 337 198 341
rect 206 338 208 341
rect 231 339 237 341
rect 162 328 164 336
rect 178 332 180 336
rect 171 330 180 332
rect 192 335 198 337
rect 192 333 194 335
rect 196 333 198 335
rect 192 331 198 333
rect 202 336 208 338
rect 202 334 204 336
rect 206 334 208 336
rect 202 332 208 334
rect 171 328 173 330
rect 175 328 180 330
rect 58 316 60 319
rect 31 310 33 315
rect 38 310 40 315
rect 58 314 63 316
rect 61 306 63 314
rect 74 310 76 314
rect 84 306 86 314
rect 122 313 124 317
rect 171 326 180 328
rect 196 328 198 331
rect 178 323 180 326
rect 188 323 190 327
rect 196 326 200 328
rect 198 323 200 326
rect 205 323 207 332
rect 235 326 237 339
rect 245 337 247 348
rect 332 368 334 372
rect 342 368 344 372
rect 349 368 351 372
rect 359 368 361 372
rect 366 368 368 372
rect 406 368 408 372
rect 416 368 418 372
rect 423 368 425 372
rect 433 368 435 372
rect 440 368 442 372
rect 480 368 482 372
rect 490 368 492 372
rect 497 368 499 372
rect 507 368 509 372
rect 514 368 516 372
rect 303 358 305 363
rect 283 344 285 347
rect 279 342 285 344
rect 255 337 257 341
rect 279 340 281 342
rect 283 340 285 342
rect 279 338 285 340
rect 241 335 247 337
rect 241 333 243 335
rect 245 333 247 335
rect 241 331 247 333
rect 251 335 257 337
rect 251 333 253 335
rect 255 333 257 335
rect 251 331 257 333
rect 242 326 244 331
rect 255 326 257 331
rect 283 328 285 338
rect 290 337 292 347
rect 379 355 385 357
rect 379 353 381 355
rect 383 353 385 355
rect 303 337 305 340
rect 289 335 295 337
rect 289 333 291 335
rect 293 333 295 335
rect 289 331 295 333
rect 299 335 305 337
rect 299 333 301 335
rect 303 333 305 335
rect 299 331 305 333
rect 332 332 334 350
rect 342 342 344 352
rect 339 340 345 342
rect 339 338 341 340
rect 343 338 345 340
rect 339 336 345 338
rect 349 337 351 352
rect 359 347 361 352
rect 356 345 362 347
rect 356 343 358 345
rect 360 343 362 345
rect 356 341 362 343
rect 366 337 368 352
rect 376 351 385 353
rect 376 348 378 351
rect 453 355 459 357
rect 453 353 455 355
rect 457 353 459 355
rect 293 328 295 331
rect 303 328 305 331
rect 331 330 337 332
rect 331 328 333 330
rect 335 328 337 330
rect 162 316 164 319
rect 94 306 96 311
rect 101 306 103 311
rect 61 304 86 306
rect 135 310 137 315
rect 142 310 144 315
rect 162 314 167 316
rect 165 306 167 314
rect 178 310 180 314
rect 188 306 190 314
rect 198 306 200 311
rect 205 306 207 311
rect 235 310 237 315
rect 242 310 244 315
rect 165 304 190 306
rect 255 313 257 317
rect 283 317 285 322
rect 293 317 295 322
rect 331 326 337 328
rect 332 323 334 326
rect 303 314 305 319
rect 342 322 344 336
rect 349 335 361 337
rect 349 329 355 331
rect 349 327 351 329
rect 353 327 355 329
rect 349 325 355 327
rect 349 322 351 325
rect 359 322 361 335
rect 366 330 372 337
rect 366 328 368 330
rect 370 328 372 330
rect 366 326 372 328
rect 366 322 368 326
rect 376 322 378 340
rect 406 332 408 350
rect 416 342 418 352
rect 413 340 419 342
rect 413 338 415 340
rect 417 338 419 340
rect 413 336 419 338
rect 423 337 425 352
rect 433 347 435 352
rect 430 345 436 347
rect 430 343 432 345
rect 434 343 436 345
rect 430 341 436 343
rect 440 337 442 352
rect 450 351 459 353
rect 450 348 452 351
rect 527 355 533 357
rect 527 353 529 355
rect 531 353 533 355
rect 405 330 411 332
rect 405 328 407 330
rect 409 328 411 330
rect 405 326 411 328
rect 406 323 408 326
rect 332 309 334 314
rect 342 309 344 314
rect 349 309 351 314
rect 359 306 361 314
rect 366 310 368 314
rect 376 306 378 316
rect 416 322 418 336
rect 423 335 435 337
rect 423 329 429 331
rect 423 327 425 329
rect 427 327 429 329
rect 423 325 429 327
rect 423 322 425 325
rect 433 322 435 335
rect 440 335 446 337
rect 440 333 442 335
rect 444 333 446 335
rect 440 331 446 333
rect 440 322 442 331
rect 450 322 452 340
rect 480 332 482 350
rect 490 342 492 352
rect 487 340 493 342
rect 487 338 489 340
rect 491 338 493 340
rect 487 336 493 338
rect 497 337 499 352
rect 507 347 509 352
rect 504 345 510 347
rect 504 343 506 345
rect 508 343 510 345
rect 504 341 510 343
rect 514 337 516 352
rect 524 351 533 353
rect 524 348 526 351
rect 479 330 485 332
rect 479 328 481 330
rect 483 328 485 330
rect 479 326 485 328
rect 480 323 482 326
rect 406 309 408 314
rect 416 309 418 314
rect 423 309 425 314
rect 359 304 378 306
rect 433 306 435 314
rect 440 310 442 314
rect 450 306 452 316
rect 490 322 492 336
rect 497 335 509 337
rect 497 329 503 331
rect 497 327 499 329
rect 501 327 503 329
rect 497 325 503 327
rect 497 322 499 325
rect 507 322 509 335
rect 514 335 520 337
rect 514 333 516 335
rect 518 333 520 335
rect 514 331 520 333
rect 514 322 516 331
rect 524 322 526 340
rect 480 309 482 314
rect 490 309 492 314
rect 497 309 499 314
rect 433 304 452 306
rect 507 306 509 314
rect 514 310 516 314
rect 524 306 526 316
rect 507 304 526 306
rect -22 285 -20 290
rect -12 282 -10 287
rect -2 282 0 287
rect 18 287 20 291
rect 31 289 33 294
rect 38 289 40 294
rect 61 298 86 300
rect 61 290 63 298
rect 74 290 76 294
rect 84 290 86 298
rect 94 293 96 298
rect 101 293 103 298
rect 58 288 63 290
rect 58 285 60 288
rect -22 273 -20 276
rect -12 273 -10 276
rect -22 271 -16 273
rect -22 269 -20 271
rect -18 269 -16 271
rect -22 267 -16 269
rect -12 271 -6 273
rect -12 269 -10 271
rect -8 269 -6 271
rect -12 267 -6 269
rect -22 264 -20 267
rect -9 257 -7 267
rect -2 266 0 276
rect 18 273 20 278
rect 31 273 33 278
rect 18 271 24 273
rect 18 269 20 271
rect 22 269 24 271
rect 18 267 24 269
rect 28 271 34 273
rect 28 269 30 271
rect 32 269 34 271
rect 28 267 34 269
rect -2 264 4 266
rect -2 262 0 264
rect 2 262 4 264
rect 18 263 20 267
rect -2 260 4 262
rect -2 257 0 260
rect -22 241 -20 246
rect 28 256 30 267
rect 38 265 40 278
rect 122 287 124 291
rect 135 289 137 294
rect 142 289 144 294
rect 165 298 190 300
rect 165 290 167 298
rect 178 290 180 294
rect 188 290 190 298
rect 198 293 200 298
rect 205 293 207 298
rect 74 278 76 281
rect 67 276 76 278
rect 84 277 86 281
rect 94 278 96 281
rect 58 268 60 276
rect 67 274 69 276
rect 71 274 76 276
rect 67 272 76 274
rect 92 276 96 278
rect 92 273 94 276
rect 74 268 76 272
rect 88 271 94 273
rect 101 272 103 281
rect 162 288 167 290
rect 162 285 164 288
rect 122 273 124 278
rect 135 273 137 278
rect 88 269 90 271
rect 92 269 94 271
rect 55 266 68 268
rect 74 266 84 268
rect 88 267 94 269
rect 55 265 57 266
rect 38 263 44 265
rect 38 261 40 263
rect 42 261 44 263
rect 38 259 44 261
rect 51 263 57 265
rect 66 263 68 266
rect 82 263 84 266
rect 92 263 94 267
rect 98 270 104 272
rect 98 268 100 270
rect 102 268 104 270
rect 98 266 104 268
rect 102 263 104 266
rect 122 271 128 273
rect 122 269 124 271
rect 126 269 128 271
rect 122 267 128 269
rect 132 271 138 273
rect 132 269 134 271
rect 136 269 138 271
rect 132 267 138 269
rect 122 263 124 267
rect 51 261 53 263
rect 55 261 57 263
rect 51 259 57 261
rect 38 256 40 259
rect 18 241 20 245
rect 28 238 30 243
rect 38 238 40 243
rect -9 232 -7 236
rect -2 232 0 236
rect 82 241 84 245
rect 92 241 94 245
rect 66 232 68 236
rect 132 256 134 267
rect 142 265 144 278
rect 235 289 237 294
rect 242 289 244 294
rect 359 298 378 300
rect 178 278 180 281
rect 171 276 180 278
rect 188 277 190 281
rect 198 278 200 281
rect 162 268 164 276
rect 171 274 173 276
rect 175 274 180 276
rect 171 272 180 274
rect 196 276 200 278
rect 196 273 198 276
rect 178 268 180 272
rect 192 271 198 273
rect 205 272 207 281
rect 255 287 257 291
rect 332 290 334 295
rect 342 290 344 295
rect 349 290 351 295
rect 359 290 361 298
rect 366 290 368 294
rect 283 282 285 287
rect 293 282 295 287
rect 303 285 305 290
rect 192 269 194 271
rect 196 269 198 271
rect 159 266 172 268
rect 178 266 188 268
rect 192 267 198 269
rect 159 265 161 266
rect 142 263 148 265
rect 142 261 144 263
rect 146 261 148 263
rect 142 259 148 261
rect 155 263 161 265
rect 170 263 172 266
rect 186 263 188 266
rect 196 263 198 267
rect 202 270 208 272
rect 202 268 204 270
rect 206 268 208 270
rect 202 266 208 268
rect 206 263 208 266
rect 235 265 237 278
rect 242 273 244 278
rect 255 273 257 278
rect 376 288 378 298
rect 433 298 452 300
rect 406 290 408 295
rect 416 290 418 295
rect 423 290 425 295
rect 433 290 435 298
rect 440 290 442 294
rect 332 278 334 281
rect 331 276 337 278
rect 241 271 247 273
rect 241 269 243 271
rect 245 269 247 271
rect 241 267 247 269
rect 251 271 257 273
rect 251 269 253 271
rect 255 269 257 271
rect 251 267 257 269
rect 231 263 237 265
rect 155 261 157 263
rect 159 261 161 263
rect 155 259 161 261
rect 142 256 144 259
rect 122 241 124 245
rect 132 238 134 243
rect 142 238 144 243
rect 102 232 104 236
rect 186 241 188 245
rect 196 241 198 245
rect 170 232 172 236
rect 231 261 233 263
rect 235 261 237 263
rect 231 259 237 261
rect 235 256 237 259
rect 245 256 247 267
rect 255 263 257 267
rect 283 266 285 276
rect 293 273 295 276
rect 303 273 305 276
rect 289 271 295 273
rect 289 269 291 271
rect 293 269 295 271
rect 289 267 295 269
rect 299 271 305 273
rect 331 274 333 276
rect 335 274 337 276
rect 331 272 337 274
rect 299 269 301 271
rect 303 269 305 271
rect 299 267 305 269
rect 279 264 285 266
rect 279 262 281 264
rect 283 262 285 264
rect 279 260 285 262
rect 283 257 285 260
rect 290 257 292 267
rect 303 264 305 267
rect 235 238 237 243
rect 245 238 247 243
rect 255 241 257 245
rect 206 232 208 236
rect 332 254 334 272
rect 342 268 344 282
rect 349 279 351 282
rect 349 277 355 279
rect 349 275 351 277
rect 353 275 355 277
rect 349 273 355 275
rect 359 269 361 282
rect 339 266 345 268
rect 339 264 341 266
rect 343 264 345 266
rect 339 262 345 264
rect 349 267 361 269
rect 366 278 368 282
rect 366 276 372 278
rect 366 274 368 276
rect 370 274 372 276
rect 366 267 372 274
rect 303 241 305 246
rect 283 232 285 236
rect 290 232 292 236
rect 342 252 344 262
rect 349 252 351 267
rect 356 261 362 263
rect 356 259 358 261
rect 360 259 362 261
rect 356 257 362 259
rect 359 252 361 257
rect 366 252 368 267
rect 376 264 378 282
rect 450 288 452 298
rect 507 298 526 300
rect 480 290 482 295
rect 490 290 492 295
rect 497 290 499 295
rect 507 290 509 298
rect 514 290 516 294
rect 406 278 408 281
rect 405 276 411 278
rect 405 274 407 276
rect 409 274 411 276
rect 405 272 411 274
rect 376 253 378 256
rect 406 254 408 272
rect 416 268 418 282
rect 423 279 425 282
rect 423 277 429 279
rect 423 275 425 277
rect 427 275 429 277
rect 423 273 429 275
rect 433 269 435 282
rect 413 266 419 268
rect 413 264 415 266
rect 417 264 419 266
rect 413 262 419 264
rect 423 267 435 269
rect 440 273 442 282
rect 440 271 446 273
rect 440 269 442 271
rect 444 269 446 271
rect 440 267 446 269
rect 376 251 385 253
rect 379 249 381 251
rect 383 249 385 251
rect 379 247 385 249
rect 416 252 418 262
rect 423 252 425 267
rect 430 261 436 263
rect 430 259 432 261
rect 434 259 436 261
rect 430 257 436 259
rect 433 252 435 257
rect 440 252 442 267
rect 450 264 452 282
rect 524 288 526 298
rect 480 278 482 281
rect 479 276 485 278
rect 479 274 481 276
rect 483 274 485 276
rect 479 272 485 274
rect 450 253 452 256
rect 480 254 482 272
rect 490 268 492 282
rect 497 279 499 282
rect 497 277 503 279
rect 497 275 499 277
rect 501 275 503 277
rect 497 273 503 275
rect 507 269 509 282
rect 487 266 493 268
rect 487 264 489 266
rect 491 264 493 266
rect 487 262 493 264
rect 497 267 509 269
rect 514 273 516 282
rect 514 271 520 273
rect 514 269 516 271
rect 518 269 520 271
rect 514 267 520 269
rect 450 251 459 253
rect 453 249 455 251
rect 457 249 459 251
rect 453 247 459 249
rect 490 252 492 262
rect 497 252 499 267
rect 504 261 510 263
rect 504 259 506 261
rect 508 259 510 261
rect 504 257 510 259
rect 507 252 509 257
rect 514 252 516 267
rect 524 264 526 282
rect 524 253 526 256
rect 524 251 533 253
rect 527 249 529 251
rect 531 249 533 251
rect 527 247 533 249
rect 332 232 334 236
rect 342 232 344 236
rect 349 232 351 236
rect 359 232 361 236
rect 366 232 368 236
rect 406 232 408 236
rect 416 232 418 236
rect 423 232 425 236
rect 433 232 435 236
rect 440 232 442 236
rect 480 232 482 236
rect 490 232 492 236
rect 497 232 499 236
rect 507 232 509 236
rect 514 232 516 236
rect -9 224 -7 228
rect -2 224 0 228
rect -22 214 -20 219
rect 66 224 68 228
rect 18 215 20 219
rect 28 217 30 222
rect 38 217 40 222
rect -22 193 -20 196
rect -9 193 -7 203
rect -2 200 0 203
rect -2 198 4 200
rect -2 196 0 198
rect 2 196 4 198
rect -2 194 4 196
rect -22 191 -16 193
rect -22 189 -20 191
rect -18 189 -16 191
rect -22 187 -16 189
rect -12 191 -6 193
rect -12 189 -10 191
rect -8 189 -6 191
rect -12 187 -6 189
rect -22 184 -20 187
rect -12 184 -10 187
rect -2 184 0 194
rect 18 193 20 197
rect 28 193 30 204
rect 38 201 40 204
rect 38 199 44 201
rect 38 197 40 199
rect 42 197 44 199
rect 38 195 44 197
rect 51 199 57 201
rect 51 197 53 199
rect 55 197 57 199
rect 102 224 104 228
rect 82 215 84 219
rect 92 215 94 219
rect 170 224 172 228
rect 122 215 124 219
rect 132 217 134 222
rect 142 217 144 222
rect 51 195 57 197
rect 18 191 24 193
rect 18 189 20 191
rect 22 189 24 191
rect 18 187 24 189
rect 28 191 34 193
rect 28 189 30 191
rect 32 189 34 191
rect 28 187 34 189
rect 18 182 20 187
rect 31 182 33 187
rect 38 182 40 195
rect 55 194 57 195
rect 66 194 68 197
rect 82 194 84 197
rect 55 192 68 194
rect 74 192 84 194
rect 92 193 94 197
rect 102 194 104 197
rect 58 184 60 192
rect 74 188 76 192
rect 67 186 76 188
rect 88 191 94 193
rect 88 189 90 191
rect 92 189 94 191
rect 88 187 94 189
rect 98 192 104 194
rect 98 190 100 192
rect 102 190 104 192
rect 98 188 104 190
rect 122 193 124 197
rect 132 193 134 204
rect 142 201 144 204
rect 142 199 148 201
rect 142 197 144 199
rect 146 197 148 199
rect 142 195 148 197
rect 155 199 161 201
rect 155 197 157 199
rect 159 197 161 199
rect 206 224 208 228
rect 186 215 188 219
rect 196 215 198 219
rect 283 224 285 228
rect 290 224 292 228
rect 235 217 237 222
rect 245 217 247 222
rect 255 215 257 219
rect 235 201 237 204
rect 231 199 237 201
rect 231 197 233 199
rect 235 197 237 199
rect 155 195 161 197
rect 122 191 128 193
rect 122 189 124 191
rect 126 189 128 191
rect 67 184 69 186
rect 71 184 76 186
rect -22 170 -20 175
rect -12 173 -10 178
rect -2 173 0 178
rect 18 169 20 173
rect 67 182 76 184
rect 92 184 94 187
rect 74 179 76 182
rect 84 179 86 183
rect 92 182 96 184
rect 94 179 96 182
rect 101 179 103 188
rect 122 187 128 189
rect 132 191 138 193
rect 132 189 134 191
rect 136 189 138 191
rect 132 187 138 189
rect 122 182 124 187
rect 135 182 137 187
rect 142 182 144 195
rect 159 194 161 195
rect 170 194 172 197
rect 186 194 188 197
rect 159 192 172 194
rect 178 192 188 194
rect 196 193 198 197
rect 206 194 208 197
rect 231 195 237 197
rect 162 184 164 192
rect 178 188 180 192
rect 171 186 180 188
rect 192 191 198 193
rect 192 189 194 191
rect 196 189 198 191
rect 192 187 198 189
rect 202 192 208 194
rect 202 190 204 192
rect 206 190 208 192
rect 202 188 208 190
rect 171 184 173 186
rect 175 184 180 186
rect 58 172 60 175
rect 31 166 33 171
rect 38 166 40 171
rect 58 170 63 172
rect 61 162 63 170
rect 74 166 76 170
rect 84 162 86 170
rect 122 169 124 173
rect 171 182 180 184
rect 196 184 198 187
rect 178 179 180 182
rect 188 179 190 183
rect 196 182 200 184
rect 198 179 200 182
rect 205 179 207 188
rect 235 182 237 195
rect 245 193 247 204
rect 332 224 334 228
rect 342 224 344 228
rect 349 224 351 228
rect 359 224 361 228
rect 366 224 368 228
rect 406 224 408 228
rect 416 224 418 228
rect 423 224 425 228
rect 433 224 435 228
rect 440 224 442 228
rect 480 224 482 228
rect 490 224 492 228
rect 497 224 499 228
rect 507 224 509 228
rect 514 224 516 228
rect 303 214 305 219
rect 283 200 285 203
rect 279 198 285 200
rect 255 193 257 197
rect 279 196 281 198
rect 283 196 285 198
rect 279 194 285 196
rect 241 191 247 193
rect 241 189 243 191
rect 245 189 247 191
rect 241 187 247 189
rect 251 191 257 193
rect 251 189 253 191
rect 255 189 257 191
rect 251 187 257 189
rect 242 182 244 187
rect 255 182 257 187
rect 283 184 285 194
rect 290 193 292 203
rect 379 211 385 213
rect 379 209 381 211
rect 383 209 385 211
rect 303 193 305 196
rect 289 191 295 193
rect 289 189 291 191
rect 293 189 295 191
rect 289 187 295 189
rect 299 191 305 193
rect 299 189 301 191
rect 303 189 305 191
rect 299 187 305 189
rect 332 188 334 206
rect 342 198 344 208
rect 339 196 345 198
rect 339 194 341 196
rect 343 194 345 196
rect 339 192 345 194
rect 349 193 351 208
rect 359 203 361 208
rect 356 201 362 203
rect 356 199 358 201
rect 360 199 362 201
rect 356 197 362 199
rect 366 193 368 208
rect 376 207 385 209
rect 376 204 378 207
rect 453 211 459 213
rect 453 209 455 211
rect 457 209 459 211
rect 293 184 295 187
rect 303 184 305 187
rect 331 186 337 188
rect 331 184 333 186
rect 335 184 337 186
rect 162 172 164 175
rect 94 162 96 167
rect 101 162 103 167
rect 61 160 86 162
rect 135 166 137 171
rect 142 166 144 171
rect 162 170 167 172
rect 165 162 167 170
rect 178 166 180 170
rect 188 162 190 170
rect 198 162 200 167
rect 205 162 207 167
rect 235 166 237 171
rect 242 166 244 171
rect 165 160 190 162
rect 255 169 257 173
rect 283 173 285 178
rect 293 173 295 178
rect 331 182 337 184
rect 332 179 334 182
rect 303 170 305 175
rect 342 178 344 192
rect 349 191 361 193
rect 349 185 355 187
rect 349 183 351 185
rect 353 183 355 185
rect 349 181 355 183
rect 349 178 351 181
rect 359 178 361 191
rect 366 186 372 193
rect 366 184 368 186
rect 370 184 372 186
rect 366 182 372 184
rect 366 178 368 182
rect 376 178 378 196
rect 406 188 408 206
rect 416 198 418 208
rect 413 196 419 198
rect 413 194 415 196
rect 417 194 419 196
rect 413 192 419 194
rect 423 193 425 208
rect 433 203 435 208
rect 430 201 436 203
rect 430 199 432 201
rect 434 199 436 201
rect 430 197 436 199
rect 440 193 442 208
rect 450 207 459 209
rect 450 204 452 207
rect 527 211 533 213
rect 527 209 529 211
rect 531 209 533 211
rect 405 186 411 188
rect 405 184 407 186
rect 409 184 411 186
rect 405 182 411 184
rect 406 179 408 182
rect 332 165 334 170
rect 342 165 344 170
rect 349 165 351 170
rect 359 162 361 170
rect 366 166 368 170
rect 376 162 378 172
rect 416 178 418 192
rect 423 191 435 193
rect 423 185 429 187
rect 423 183 425 185
rect 427 183 429 185
rect 423 181 429 183
rect 423 178 425 181
rect 433 178 435 191
rect 440 191 446 193
rect 440 189 442 191
rect 444 189 446 191
rect 440 187 446 189
rect 440 178 442 187
rect 450 178 452 196
rect 480 188 482 206
rect 490 198 492 208
rect 487 196 493 198
rect 487 194 489 196
rect 491 194 493 196
rect 487 192 493 194
rect 497 193 499 208
rect 507 203 509 208
rect 504 201 510 203
rect 504 199 506 201
rect 508 199 510 201
rect 504 197 510 199
rect 514 193 516 208
rect 524 207 533 209
rect 524 204 526 207
rect 479 186 485 188
rect 479 184 481 186
rect 483 184 485 186
rect 479 182 485 184
rect 480 179 482 182
rect 406 165 408 170
rect 416 165 418 170
rect 423 165 425 170
rect 359 160 378 162
rect 433 162 435 170
rect 440 166 442 170
rect 450 162 452 172
rect 490 178 492 192
rect 497 191 509 193
rect 497 185 503 187
rect 497 183 499 185
rect 501 183 503 185
rect 497 181 503 183
rect 497 178 499 181
rect 507 178 509 191
rect 514 191 520 193
rect 514 189 516 191
rect 518 189 520 191
rect 514 187 520 189
rect 514 178 516 187
rect 524 178 526 196
rect 480 165 482 170
rect 490 165 492 170
rect 497 165 499 170
rect 433 160 452 162
rect 507 162 509 170
rect 514 166 516 170
rect 524 162 526 172
rect 507 160 526 162
<< ndif >>
rect -18 437 -12 439
rect -18 435 -16 437
rect -14 435 -12 437
rect -18 433 -12 435
rect 1 437 7 439
rect 22 441 29 443
rect 22 439 24 441
rect 26 439 29 441
rect 1 435 3 437
rect 5 435 7 437
rect 1 433 7 435
rect -18 429 -14 433
rect -27 426 -22 429
rect -29 424 -22 426
rect -29 422 -27 424
rect -25 422 -22 424
rect -29 420 -22 422
rect -20 426 -14 429
rect 2 426 7 433
rect 22 433 29 439
rect 105 441 111 443
rect 105 439 107 441
rect 109 439 111 441
rect 105 437 111 439
rect 126 441 133 443
rect 126 439 128 441
rect 130 439 133 441
rect 89 434 94 437
rect 22 431 31 433
rect -20 420 -12 426
rect -10 424 -2 426
rect -10 422 -7 424
rect -5 422 -2 424
rect -10 420 -2 422
rect 0 420 7 426
rect 11 429 18 431
rect 11 427 13 429
rect 15 427 18 429
rect 11 425 18 427
rect 13 422 18 425
rect 20 422 31 431
rect 33 422 38 433
rect 40 431 47 433
rect 40 429 43 431
rect 45 429 47 431
rect 65 432 74 434
rect 65 430 67 432
rect 69 430 74 432
rect 65 429 74 430
rect 40 427 47 429
rect 40 422 45 427
rect 53 426 58 429
rect 51 424 58 426
rect 51 422 53 424
rect 55 422 58 424
rect 51 420 58 422
rect 60 425 74 429
rect 76 429 84 434
rect 76 427 79 429
rect 81 427 84 429
rect 76 425 84 427
rect 86 431 94 434
rect 86 429 89 431
rect 91 429 94 431
rect 86 425 94 429
rect 96 425 101 437
rect 103 425 111 437
rect 126 433 133 439
rect 209 441 215 443
rect 209 439 211 441
rect 213 439 215 441
rect 209 437 215 439
rect 246 441 253 443
rect 246 439 249 441
rect 251 439 253 441
rect 193 434 198 437
rect 126 431 135 433
rect 115 429 122 431
rect 115 427 117 429
rect 119 427 122 429
rect 115 425 122 427
rect 60 420 65 425
rect 117 422 122 425
rect 124 422 135 431
rect 137 422 142 433
rect 144 431 151 433
rect 144 429 147 431
rect 149 429 151 431
rect 169 432 178 434
rect 169 430 171 432
rect 173 430 178 432
rect 169 429 178 430
rect 144 427 151 429
rect 144 422 149 427
rect 157 426 162 429
rect 155 424 162 426
rect 155 422 157 424
rect 159 422 162 424
rect 155 420 162 422
rect 164 425 178 429
rect 180 429 188 434
rect 180 427 183 429
rect 185 427 188 429
rect 180 425 188 427
rect 190 431 198 434
rect 190 429 193 431
rect 195 429 198 431
rect 190 425 198 429
rect 200 425 205 437
rect 207 425 215 437
rect 246 433 253 439
rect 276 437 282 439
rect 276 435 278 437
rect 280 435 282 437
rect 228 431 235 433
rect 228 429 230 431
rect 232 429 235 431
rect 228 427 235 429
rect 164 420 169 425
rect 230 422 235 427
rect 237 422 242 433
rect 244 431 253 433
rect 276 433 282 435
rect 295 437 301 439
rect 295 435 297 437
rect 299 435 301 437
rect 295 433 301 435
rect 244 422 255 431
rect 257 429 264 431
rect 257 427 260 429
rect 262 427 264 429
rect 257 425 264 427
rect 276 426 281 433
rect 297 429 301 433
rect 327 431 332 434
rect 325 429 332 431
rect 297 426 303 429
rect 257 422 262 425
rect 276 420 283 426
rect 285 424 293 426
rect 285 422 288 424
rect 290 422 293 424
rect 285 420 293 422
rect 295 420 303 426
rect 305 426 310 429
rect 325 427 327 429
rect 329 427 332 429
rect 305 424 312 426
rect 325 425 332 427
rect 334 432 342 434
rect 334 430 337 432
rect 339 430 342 432
rect 334 426 342 430
rect 344 426 349 434
rect 351 432 359 434
rect 351 430 354 432
rect 356 430 359 432
rect 351 426 359 430
rect 361 426 366 434
rect 368 432 374 434
rect 368 430 376 432
rect 368 428 371 430
rect 373 428 376 430
rect 368 426 376 428
rect 378 430 385 432
rect 401 431 406 434
rect 378 428 381 430
rect 383 428 385 430
rect 378 426 385 428
rect 399 429 406 431
rect 399 427 401 429
rect 403 427 406 429
rect 334 425 339 426
rect 305 422 308 424
rect 310 422 312 424
rect 305 420 312 422
rect 399 425 406 427
rect 408 432 416 434
rect 408 430 411 432
rect 413 430 416 432
rect 408 426 416 430
rect 418 426 423 434
rect 425 432 433 434
rect 425 430 428 432
rect 430 430 433 432
rect 425 426 433 430
rect 435 426 440 434
rect 442 432 448 434
rect 442 430 450 432
rect 442 428 445 430
rect 447 428 450 430
rect 442 426 450 428
rect 452 430 459 432
rect 475 431 480 434
rect 452 428 455 430
rect 457 428 459 430
rect 452 426 459 428
rect 473 429 480 431
rect 473 427 475 429
rect 477 427 480 429
rect 408 425 413 426
rect 473 425 480 427
rect 482 432 490 434
rect 482 430 485 432
rect 487 430 490 432
rect 482 426 490 430
rect 492 426 497 434
rect 499 432 507 434
rect 499 430 502 432
rect 504 430 507 432
rect 499 426 507 430
rect 509 426 514 434
rect 516 432 522 434
rect 516 430 524 432
rect 516 428 519 430
rect 521 428 524 430
rect 516 426 524 428
rect 526 430 533 432
rect 526 428 529 430
rect 531 428 533 430
rect 526 426 533 428
rect 482 425 487 426
rect -29 326 -22 328
rect -29 324 -27 326
rect -25 324 -22 326
rect -29 322 -22 324
rect -27 319 -22 322
rect -20 322 -12 328
rect -10 326 -2 328
rect -10 324 -7 326
rect -5 324 -2 326
rect -10 322 -2 324
rect 0 322 7 328
rect 51 326 58 328
rect 13 323 18 326
rect -20 319 -14 322
rect -18 315 -14 319
rect 2 315 7 322
rect 11 321 18 323
rect 11 319 13 321
rect 15 319 18 321
rect 11 317 18 319
rect 20 317 31 326
rect -18 313 -12 315
rect -18 311 -16 313
rect -14 311 -12 313
rect -18 309 -12 311
rect 1 313 7 315
rect 22 315 31 317
rect 33 315 38 326
rect 40 321 45 326
rect 51 324 53 326
rect 55 324 58 326
rect 51 322 58 324
rect 40 319 47 321
rect 53 319 58 322
rect 60 323 65 328
rect 155 326 162 328
rect 117 323 122 326
rect 60 319 74 323
rect 40 317 43 319
rect 45 317 47 319
rect 40 315 47 317
rect 65 318 74 319
rect 65 316 67 318
rect 69 316 74 318
rect 1 311 3 313
rect 5 311 7 313
rect 1 309 7 311
rect 22 309 29 315
rect 65 314 74 316
rect 76 321 84 323
rect 76 319 79 321
rect 81 319 84 321
rect 76 314 84 319
rect 86 319 94 323
rect 86 317 89 319
rect 91 317 94 319
rect 86 314 94 317
rect 22 307 24 309
rect 26 307 29 309
rect 22 305 29 307
rect 89 311 94 314
rect 96 311 101 323
rect 103 311 111 323
rect 115 321 122 323
rect 115 319 117 321
rect 119 319 122 321
rect 115 317 122 319
rect 124 317 135 326
rect 126 315 135 317
rect 137 315 142 326
rect 144 321 149 326
rect 155 324 157 326
rect 159 324 162 326
rect 155 322 162 324
rect 144 319 151 321
rect 157 319 162 322
rect 164 323 169 328
rect 164 319 178 323
rect 144 317 147 319
rect 149 317 151 319
rect 144 315 151 317
rect 169 318 178 319
rect 169 316 171 318
rect 173 316 178 318
rect 105 309 111 311
rect 105 307 107 309
rect 109 307 111 309
rect 105 305 111 307
rect 126 309 133 315
rect 169 314 178 316
rect 180 321 188 323
rect 180 319 183 321
rect 185 319 188 321
rect 180 314 188 319
rect 190 319 198 323
rect 190 317 193 319
rect 195 317 198 319
rect 190 314 198 317
rect 126 307 128 309
rect 130 307 133 309
rect 126 305 133 307
rect 193 311 198 314
rect 200 311 205 323
rect 207 311 215 323
rect 230 321 235 326
rect 228 319 235 321
rect 228 317 230 319
rect 232 317 235 319
rect 228 315 235 317
rect 237 315 242 326
rect 244 317 255 326
rect 257 323 262 326
rect 257 321 264 323
rect 257 319 260 321
rect 262 319 264 321
rect 257 317 264 319
rect 276 322 283 328
rect 285 326 293 328
rect 285 324 288 326
rect 290 324 293 326
rect 285 322 293 324
rect 295 322 303 328
rect 244 315 253 317
rect 209 309 215 311
rect 209 307 211 309
rect 213 307 215 309
rect 209 305 215 307
rect 246 309 253 315
rect 276 315 281 322
rect 297 319 303 322
rect 305 326 312 328
rect 305 324 308 326
rect 310 324 312 326
rect 305 322 312 324
rect 305 319 310 322
rect 325 321 332 323
rect 325 319 327 321
rect 329 319 332 321
rect 297 315 301 319
rect 276 313 282 315
rect 276 311 278 313
rect 280 311 282 313
rect 246 307 249 309
rect 251 307 253 309
rect 246 305 253 307
rect 276 309 282 311
rect 295 313 301 315
rect 325 317 332 319
rect 327 314 332 317
rect 334 322 339 323
rect 334 318 342 322
rect 334 316 337 318
rect 339 316 342 318
rect 334 314 342 316
rect 344 314 349 322
rect 351 318 359 322
rect 351 316 354 318
rect 356 316 359 318
rect 351 314 359 316
rect 361 314 366 322
rect 368 320 376 322
rect 368 318 371 320
rect 373 318 376 320
rect 368 316 376 318
rect 378 320 385 322
rect 378 318 381 320
rect 383 318 385 320
rect 378 316 385 318
rect 399 321 406 323
rect 399 319 401 321
rect 403 319 406 321
rect 399 317 406 319
rect 368 314 374 316
rect 295 311 297 313
rect 299 311 301 313
rect 295 309 301 311
rect 401 314 406 317
rect 408 322 413 323
rect 408 318 416 322
rect 408 316 411 318
rect 413 316 416 318
rect 408 314 416 316
rect 418 314 423 322
rect 425 318 433 322
rect 425 316 428 318
rect 430 316 433 318
rect 425 314 433 316
rect 435 314 440 322
rect 442 320 450 322
rect 442 318 445 320
rect 447 318 450 320
rect 442 316 450 318
rect 452 320 459 322
rect 452 318 455 320
rect 457 318 459 320
rect 452 316 459 318
rect 473 321 480 323
rect 473 319 475 321
rect 477 319 480 321
rect 473 317 480 319
rect 442 314 448 316
rect 475 314 480 317
rect 482 322 487 323
rect 482 318 490 322
rect 482 316 485 318
rect 487 316 490 318
rect 482 314 490 316
rect 492 314 497 322
rect 499 318 507 322
rect 499 316 502 318
rect 504 316 507 318
rect 499 314 507 316
rect 509 314 514 322
rect 516 320 524 322
rect 516 318 519 320
rect 521 318 524 320
rect 516 316 524 318
rect 526 320 533 322
rect 526 318 529 320
rect 531 318 533 320
rect 526 316 533 318
rect 516 314 522 316
rect -18 293 -12 295
rect -18 291 -16 293
rect -14 291 -12 293
rect -18 289 -12 291
rect 1 293 7 295
rect 22 297 29 299
rect 22 295 24 297
rect 26 295 29 297
rect 1 291 3 293
rect 5 291 7 293
rect 1 289 7 291
rect -18 285 -14 289
rect -27 282 -22 285
rect -29 280 -22 282
rect -29 278 -27 280
rect -25 278 -22 280
rect -29 276 -22 278
rect -20 282 -14 285
rect 2 282 7 289
rect 22 289 29 295
rect 105 297 111 299
rect 105 295 107 297
rect 109 295 111 297
rect 105 293 111 295
rect 126 297 133 299
rect 126 295 128 297
rect 130 295 133 297
rect 89 290 94 293
rect 22 287 31 289
rect -20 276 -12 282
rect -10 280 -2 282
rect -10 278 -7 280
rect -5 278 -2 280
rect -10 276 -2 278
rect 0 276 7 282
rect 11 285 18 287
rect 11 283 13 285
rect 15 283 18 285
rect 11 281 18 283
rect 13 278 18 281
rect 20 278 31 287
rect 33 278 38 289
rect 40 287 47 289
rect 40 285 43 287
rect 45 285 47 287
rect 65 288 74 290
rect 65 286 67 288
rect 69 286 74 288
rect 65 285 74 286
rect 40 283 47 285
rect 40 278 45 283
rect 53 282 58 285
rect 51 280 58 282
rect 51 278 53 280
rect 55 278 58 280
rect 51 276 58 278
rect 60 281 74 285
rect 76 285 84 290
rect 76 283 79 285
rect 81 283 84 285
rect 76 281 84 283
rect 86 287 94 290
rect 86 285 89 287
rect 91 285 94 287
rect 86 281 94 285
rect 96 281 101 293
rect 103 281 111 293
rect 126 289 133 295
rect 209 297 215 299
rect 209 295 211 297
rect 213 295 215 297
rect 209 293 215 295
rect 246 297 253 299
rect 246 295 249 297
rect 251 295 253 297
rect 193 290 198 293
rect 126 287 135 289
rect 115 285 122 287
rect 115 283 117 285
rect 119 283 122 285
rect 115 281 122 283
rect 60 276 65 281
rect 117 278 122 281
rect 124 278 135 287
rect 137 278 142 289
rect 144 287 151 289
rect 144 285 147 287
rect 149 285 151 287
rect 169 288 178 290
rect 169 286 171 288
rect 173 286 178 288
rect 169 285 178 286
rect 144 283 151 285
rect 144 278 149 283
rect 157 282 162 285
rect 155 280 162 282
rect 155 278 157 280
rect 159 278 162 280
rect 155 276 162 278
rect 164 281 178 285
rect 180 285 188 290
rect 180 283 183 285
rect 185 283 188 285
rect 180 281 188 283
rect 190 287 198 290
rect 190 285 193 287
rect 195 285 198 287
rect 190 281 198 285
rect 200 281 205 293
rect 207 281 215 293
rect 246 289 253 295
rect 276 293 282 295
rect 276 291 278 293
rect 280 291 282 293
rect 228 287 235 289
rect 228 285 230 287
rect 232 285 235 287
rect 228 283 235 285
rect 164 276 169 281
rect 230 278 235 283
rect 237 278 242 289
rect 244 287 253 289
rect 276 289 282 291
rect 295 293 301 295
rect 295 291 297 293
rect 299 291 301 293
rect 295 289 301 291
rect 244 278 255 287
rect 257 285 264 287
rect 257 283 260 285
rect 262 283 264 285
rect 257 281 264 283
rect 276 282 281 289
rect 297 285 301 289
rect 327 287 332 290
rect 325 285 332 287
rect 297 282 303 285
rect 257 278 262 281
rect 276 276 283 282
rect 285 280 293 282
rect 285 278 288 280
rect 290 278 293 280
rect 285 276 293 278
rect 295 276 303 282
rect 305 282 310 285
rect 325 283 327 285
rect 329 283 332 285
rect 305 280 312 282
rect 325 281 332 283
rect 334 288 342 290
rect 334 286 337 288
rect 339 286 342 288
rect 334 282 342 286
rect 344 282 349 290
rect 351 288 359 290
rect 351 286 354 288
rect 356 286 359 288
rect 351 282 359 286
rect 361 282 366 290
rect 368 288 374 290
rect 368 286 376 288
rect 368 284 371 286
rect 373 284 376 286
rect 368 282 376 284
rect 378 286 385 288
rect 401 287 406 290
rect 378 284 381 286
rect 383 284 385 286
rect 378 282 385 284
rect 399 285 406 287
rect 399 283 401 285
rect 403 283 406 285
rect 334 281 339 282
rect 305 278 308 280
rect 310 278 312 280
rect 305 276 312 278
rect 399 281 406 283
rect 408 288 416 290
rect 408 286 411 288
rect 413 286 416 288
rect 408 282 416 286
rect 418 282 423 290
rect 425 288 433 290
rect 425 286 428 288
rect 430 286 433 288
rect 425 282 433 286
rect 435 282 440 290
rect 442 288 448 290
rect 442 286 450 288
rect 442 284 445 286
rect 447 284 450 286
rect 442 282 450 284
rect 452 286 459 288
rect 475 287 480 290
rect 452 284 455 286
rect 457 284 459 286
rect 452 282 459 284
rect 473 285 480 287
rect 473 283 475 285
rect 477 283 480 285
rect 408 281 413 282
rect 473 281 480 283
rect 482 288 490 290
rect 482 286 485 288
rect 487 286 490 288
rect 482 282 490 286
rect 492 282 497 290
rect 499 288 507 290
rect 499 286 502 288
rect 504 286 507 288
rect 499 282 507 286
rect 509 282 514 290
rect 516 288 522 290
rect 516 286 524 288
rect 516 284 519 286
rect 521 284 524 286
rect 516 282 524 284
rect 526 286 533 288
rect 526 284 529 286
rect 531 284 533 286
rect 526 282 533 284
rect 482 281 487 282
rect -29 182 -22 184
rect -29 180 -27 182
rect -25 180 -22 182
rect -29 178 -22 180
rect -27 175 -22 178
rect -20 178 -12 184
rect -10 182 -2 184
rect -10 180 -7 182
rect -5 180 -2 182
rect -10 178 -2 180
rect 0 178 7 184
rect 51 182 58 184
rect 13 179 18 182
rect -20 175 -14 178
rect -18 171 -14 175
rect 2 171 7 178
rect 11 177 18 179
rect 11 175 13 177
rect 15 175 18 177
rect 11 173 18 175
rect 20 173 31 182
rect -18 169 -12 171
rect -18 167 -16 169
rect -14 167 -12 169
rect -18 165 -12 167
rect 1 169 7 171
rect 22 171 31 173
rect 33 171 38 182
rect 40 177 45 182
rect 51 180 53 182
rect 55 180 58 182
rect 51 178 58 180
rect 40 175 47 177
rect 53 175 58 178
rect 60 179 65 184
rect 155 182 162 184
rect 117 179 122 182
rect 60 175 74 179
rect 40 173 43 175
rect 45 173 47 175
rect 40 171 47 173
rect 65 174 74 175
rect 65 172 67 174
rect 69 172 74 174
rect 1 167 3 169
rect 5 167 7 169
rect 1 165 7 167
rect 22 165 29 171
rect 65 170 74 172
rect 76 177 84 179
rect 76 175 79 177
rect 81 175 84 177
rect 76 170 84 175
rect 86 175 94 179
rect 86 173 89 175
rect 91 173 94 175
rect 86 170 94 173
rect 22 163 24 165
rect 26 163 29 165
rect 22 161 29 163
rect 89 167 94 170
rect 96 167 101 179
rect 103 167 111 179
rect 115 177 122 179
rect 115 175 117 177
rect 119 175 122 177
rect 115 173 122 175
rect 124 173 135 182
rect 126 171 135 173
rect 137 171 142 182
rect 144 177 149 182
rect 155 180 157 182
rect 159 180 162 182
rect 155 178 162 180
rect 144 175 151 177
rect 157 175 162 178
rect 164 179 169 184
rect 164 175 178 179
rect 144 173 147 175
rect 149 173 151 175
rect 144 171 151 173
rect 169 174 178 175
rect 169 172 171 174
rect 173 172 178 174
rect 105 165 111 167
rect 105 163 107 165
rect 109 163 111 165
rect 105 161 111 163
rect 126 165 133 171
rect 169 170 178 172
rect 180 177 188 179
rect 180 175 183 177
rect 185 175 188 177
rect 180 170 188 175
rect 190 175 198 179
rect 190 173 193 175
rect 195 173 198 175
rect 190 170 198 173
rect 126 163 128 165
rect 130 163 133 165
rect 126 161 133 163
rect 193 167 198 170
rect 200 167 205 179
rect 207 167 215 179
rect 230 177 235 182
rect 228 175 235 177
rect 228 173 230 175
rect 232 173 235 175
rect 228 171 235 173
rect 237 171 242 182
rect 244 173 255 182
rect 257 179 262 182
rect 257 177 264 179
rect 257 175 260 177
rect 262 175 264 177
rect 257 173 264 175
rect 276 178 283 184
rect 285 182 293 184
rect 285 180 288 182
rect 290 180 293 182
rect 285 178 293 180
rect 295 178 303 184
rect 244 171 253 173
rect 209 165 215 167
rect 209 163 211 165
rect 213 163 215 165
rect 209 161 215 163
rect 246 165 253 171
rect 276 171 281 178
rect 297 175 303 178
rect 305 182 312 184
rect 305 180 308 182
rect 310 180 312 182
rect 305 178 312 180
rect 305 175 310 178
rect 325 177 332 179
rect 325 175 327 177
rect 329 175 332 177
rect 297 171 301 175
rect 276 169 282 171
rect 276 167 278 169
rect 280 167 282 169
rect 246 163 249 165
rect 251 163 253 165
rect 246 161 253 163
rect 276 165 282 167
rect 295 169 301 171
rect 325 173 332 175
rect 327 170 332 173
rect 334 178 339 179
rect 334 174 342 178
rect 334 172 337 174
rect 339 172 342 174
rect 334 170 342 172
rect 344 170 349 178
rect 351 174 359 178
rect 351 172 354 174
rect 356 172 359 174
rect 351 170 359 172
rect 361 170 366 178
rect 368 176 376 178
rect 368 174 371 176
rect 373 174 376 176
rect 368 172 376 174
rect 378 176 385 178
rect 378 174 381 176
rect 383 174 385 176
rect 378 172 385 174
rect 399 177 406 179
rect 399 175 401 177
rect 403 175 406 177
rect 399 173 406 175
rect 368 170 374 172
rect 295 167 297 169
rect 299 167 301 169
rect 295 165 301 167
rect 401 170 406 173
rect 408 178 413 179
rect 408 174 416 178
rect 408 172 411 174
rect 413 172 416 174
rect 408 170 416 172
rect 418 170 423 178
rect 425 174 433 178
rect 425 172 428 174
rect 430 172 433 174
rect 425 170 433 172
rect 435 170 440 178
rect 442 176 450 178
rect 442 174 445 176
rect 447 174 450 176
rect 442 172 450 174
rect 452 176 459 178
rect 452 174 455 176
rect 457 174 459 176
rect 452 172 459 174
rect 473 177 480 179
rect 473 175 475 177
rect 477 175 480 177
rect 473 173 480 175
rect 442 170 448 172
rect 475 170 480 173
rect 482 178 487 179
rect 482 174 490 178
rect 482 172 485 174
rect 487 172 490 174
rect 482 170 490 172
rect 492 170 497 178
rect 499 174 507 178
rect 499 172 502 174
rect 504 172 507 174
rect 499 170 507 172
rect 509 170 514 178
rect 516 176 524 178
rect 516 174 519 176
rect 521 174 524 176
rect 516 172 524 174
rect 526 176 533 178
rect 526 174 529 176
rect 531 174 533 176
rect 526 172 533 174
rect 516 170 522 172
<< pdif >>
rect -27 403 -22 408
rect -29 401 -22 403
rect -29 399 -27 401
rect -25 399 -22 401
rect -29 394 -22 399
rect -29 392 -27 394
rect -25 392 -22 394
rect -29 390 -22 392
rect -20 401 -12 408
rect 11 405 18 407
rect 11 403 13 405
rect 15 403 18 405
rect -20 390 -9 401
rect -18 384 -9 390
rect -18 382 -16 384
rect -14 382 -9 384
rect -18 380 -9 382
rect -7 380 -2 401
rect 0 393 5 401
rect 11 398 18 403
rect 11 396 13 398
rect 15 396 18 398
rect 11 394 18 396
rect 0 391 7 393
rect 0 389 3 391
rect 5 389 7 391
rect 13 389 18 394
rect 20 400 26 407
rect 59 405 66 407
rect 59 403 61 405
rect 63 403 66 405
rect 59 401 66 403
rect 20 393 28 400
rect 20 391 23 393
rect 25 391 28 393
rect 20 389 28 391
rect 0 387 7 389
rect 0 380 5 387
rect 22 387 28 389
rect 30 398 38 400
rect 30 396 33 398
rect 35 396 38 398
rect 30 391 38 396
rect 30 389 33 391
rect 35 389 38 391
rect 30 387 38 389
rect 40 391 47 400
rect 40 389 43 391
rect 45 389 47 391
rect 40 387 47 389
rect 61 380 66 401
rect 68 391 82 407
rect 68 389 71 391
rect 73 389 82 391
rect 84 405 92 407
rect 84 403 87 405
rect 89 403 92 405
rect 84 398 92 403
rect 84 396 87 398
rect 89 396 92 398
rect 84 389 92 396
rect 94 398 102 407
rect 94 396 97 398
rect 99 396 102 398
rect 94 389 102 396
rect 68 384 80 389
rect 68 382 71 384
rect 73 382 80 384
rect 68 380 80 382
rect 97 380 102 389
rect 104 392 109 407
rect 115 405 122 407
rect 115 403 117 405
rect 119 403 122 405
rect 115 398 122 403
rect 115 396 117 398
rect 119 396 122 398
rect 115 394 122 396
rect 104 390 111 392
rect 104 388 107 390
rect 109 388 111 390
rect 117 389 122 394
rect 124 400 130 407
rect 163 405 170 407
rect 163 403 165 405
rect 167 403 170 405
rect 163 401 170 403
rect 124 393 132 400
rect 124 391 127 393
rect 129 391 132 393
rect 124 389 132 391
rect 104 386 111 388
rect 104 380 109 386
rect 126 387 132 389
rect 134 398 142 400
rect 134 396 137 398
rect 139 396 142 398
rect 134 391 142 396
rect 134 389 137 391
rect 139 389 142 391
rect 134 387 142 389
rect 144 391 151 400
rect 144 389 147 391
rect 149 389 151 391
rect 144 387 151 389
rect 165 380 170 401
rect 172 391 186 407
rect 172 389 175 391
rect 177 389 186 391
rect 188 405 196 407
rect 188 403 191 405
rect 193 403 196 405
rect 188 398 196 403
rect 188 396 191 398
rect 193 396 196 398
rect 188 389 196 396
rect 198 398 206 407
rect 198 396 201 398
rect 203 396 206 398
rect 198 389 206 396
rect 172 384 184 389
rect 172 382 175 384
rect 177 382 184 384
rect 172 380 184 382
rect 201 380 206 389
rect 208 392 213 407
rect 249 400 255 407
rect 208 390 215 392
rect 208 388 211 390
rect 213 388 215 390
rect 208 386 215 388
rect 228 391 235 400
rect 228 389 230 391
rect 232 389 235 391
rect 228 387 235 389
rect 237 398 245 400
rect 237 396 240 398
rect 242 396 245 398
rect 237 391 245 396
rect 237 389 240 391
rect 242 389 245 391
rect 237 387 245 389
rect 247 393 255 400
rect 247 391 250 393
rect 252 391 255 393
rect 247 389 255 391
rect 257 405 264 407
rect 257 403 260 405
rect 262 403 264 405
rect 257 398 264 403
rect 295 401 303 408
rect 257 396 260 398
rect 262 396 264 398
rect 257 394 264 396
rect 257 389 262 394
rect 278 393 283 401
rect 276 391 283 393
rect 276 389 278 391
rect 280 389 283 391
rect 247 387 253 389
rect 208 380 213 386
rect 276 387 283 389
rect 278 380 283 387
rect 285 380 290 401
rect 292 390 303 401
rect 305 403 310 408
rect 305 401 312 403
rect 305 399 308 401
rect 310 399 312 401
rect 305 394 312 399
rect 305 392 308 394
rect 310 392 312 394
rect 327 393 332 398
rect 305 390 312 392
rect 325 391 332 393
rect 292 384 301 390
rect 325 389 327 391
rect 329 389 332 391
rect 325 387 332 389
rect 292 382 297 384
rect 299 382 301 384
rect 292 380 301 382
rect 327 380 332 387
rect 334 396 339 398
rect 370 400 376 408
rect 378 406 385 408
rect 378 404 381 406
rect 383 404 385 406
rect 378 402 385 404
rect 378 400 383 402
rect 370 396 374 400
rect 334 384 342 396
rect 334 382 337 384
rect 339 382 342 384
rect 334 380 342 382
rect 344 380 349 396
rect 351 394 359 396
rect 351 392 354 394
rect 356 392 359 394
rect 351 380 359 392
rect 361 380 366 396
rect 368 392 374 396
rect 401 393 406 398
rect 368 384 375 392
rect 399 391 406 393
rect 399 389 401 391
rect 403 389 406 391
rect 399 387 406 389
rect 368 382 371 384
rect 373 382 375 384
rect 368 380 375 382
rect 401 380 406 387
rect 408 396 413 398
rect 444 400 450 408
rect 452 406 459 408
rect 452 404 455 406
rect 457 404 459 406
rect 452 402 459 404
rect 452 400 457 402
rect 444 396 448 400
rect 408 384 416 396
rect 408 382 411 384
rect 413 382 416 384
rect 408 380 416 382
rect 418 380 423 396
rect 425 394 433 396
rect 425 392 428 394
rect 430 392 433 394
rect 425 380 433 392
rect 435 380 440 396
rect 442 392 448 396
rect 475 393 480 398
rect 442 384 449 392
rect 473 391 480 393
rect 473 389 475 391
rect 477 389 480 391
rect 473 387 480 389
rect 442 382 445 384
rect 447 382 449 384
rect 442 380 449 382
rect 475 380 480 387
rect 482 396 487 398
rect 518 400 524 408
rect 526 406 533 408
rect 526 404 529 406
rect 531 404 533 406
rect 526 402 533 404
rect 526 400 531 402
rect 518 396 522 400
rect 482 384 490 396
rect 482 382 485 384
rect 487 382 490 384
rect 482 380 490 382
rect 492 380 497 396
rect 499 394 507 396
rect 499 392 502 394
rect 504 392 507 394
rect 499 380 507 392
rect 509 380 514 396
rect 516 392 522 396
rect 516 384 523 392
rect 516 382 519 384
rect 521 382 523 384
rect 516 380 523 382
rect -18 366 -9 368
rect -18 364 -16 366
rect -14 364 -9 366
rect -18 358 -9 364
rect -29 356 -22 358
rect -29 354 -27 356
rect -25 354 -22 356
rect -29 349 -22 354
rect -29 347 -27 349
rect -25 347 -22 349
rect -29 345 -22 347
rect -27 340 -22 345
rect -20 347 -9 358
rect -7 347 -2 368
rect 0 361 5 368
rect 0 359 7 361
rect 22 359 28 361
rect 0 357 3 359
rect 5 357 7 359
rect 0 355 7 357
rect 0 347 5 355
rect 13 354 18 359
rect 11 352 18 354
rect 11 350 13 352
rect 15 350 18 352
rect -20 340 -12 347
rect 11 345 18 350
rect 11 343 13 345
rect 15 343 18 345
rect 11 341 18 343
rect 20 357 28 359
rect 20 355 23 357
rect 25 355 28 357
rect 20 348 28 355
rect 30 359 38 361
rect 30 357 33 359
rect 35 357 38 359
rect 30 352 38 357
rect 30 350 33 352
rect 35 350 38 352
rect 30 348 38 350
rect 40 359 47 361
rect 40 357 43 359
rect 45 357 47 359
rect 40 348 47 357
rect 20 341 26 348
rect 61 347 66 368
rect 59 345 66 347
rect 59 343 61 345
rect 63 343 66 345
rect 59 341 66 343
rect 68 366 80 368
rect 68 364 71 366
rect 73 364 80 366
rect 68 359 80 364
rect 97 359 102 368
rect 68 357 71 359
rect 73 357 82 359
rect 68 341 82 357
rect 84 352 92 359
rect 84 350 87 352
rect 89 350 92 352
rect 84 345 92 350
rect 84 343 87 345
rect 89 343 92 345
rect 84 341 92 343
rect 94 352 102 359
rect 94 350 97 352
rect 99 350 102 352
rect 94 341 102 350
rect 104 362 109 368
rect 104 360 111 362
rect 104 358 107 360
rect 109 358 111 360
rect 126 359 132 361
rect 104 356 111 358
rect 104 341 109 356
rect 117 354 122 359
rect 115 352 122 354
rect 115 350 117 352
rect 119 350 122 352
rect 115 345 122 350
rect 115 343 117 345
rect 119 343 122 345
rect 115 341 122 343
rect 124 357 132 359
rect 124 355 127 357
rect 129 355 132 357
rect 124 348 132 355
rect 134 359 142 361
rect 134 357 137 359
rect 139 357 142 359
rect 134 352 142 357
rect 134 350 137 352
rect 139 350 142 352
rect 134 348 142 350
rect 144 359 151 361
rect 144 357 147 359
rect 149 357 151 359
rect 144 348 151 357
rect 124 341 130 348
rect 165 347 170 368
rect 163 345 170 347
rect 163 343 165 345
rect 167 343 170 345
rect 163 341 170 343
rect 172 366 184 368
rect 172 364 175 366
rect 177 364 184 366
rect 172 359 184 364
rect 201 359 206 368
rect 172 357 175 359
rect 177 357 186 359
rect 172 341 186 357
rect 188 352 196 359
rect 188 350 191 352
rect 193 350 196 352
rect 188 345 196 350
rect 188 343 191 345
rect 193 343 196 345
rect 188 341 196 343
rect 198 352 206 359
rect 198 350 201 352
rect 203 350 206 352
rect 198 341 206 350
rect 208 362 213 368
rect 208 360 215 362
rect 208 358 211 360
rect 213 358 215 360
rect 208 356 215 358
rect 228 359 235 361
rect 228 357 230 359
rect 232 357 235 359
rect 208 341 213 356
rect 228 348 235 357
rect 237 359 245 361
rect 237 357 240 359
rect 242 357 245 359
rect 237 352 245 357
rect 237 350 240 352
rect 242 350 245 352
rect 237 348 245 350
rect 247 359 253 361
rect 278 361 283 368
rect 276 359 283 361
rect 247 357 255 359
rect 247 355 250 357
rect 252 355 255 357
rect 247 348 255 355
rect 249 341 255 348
rect 257 354 262 359
rect 276 357 278 359
rect 280 357 283 359
rect 276 355 283 357
rect 257 352 264 354
rect 257 350 260 352
rect 262 350 264 352
rect 257 345 264 350
rect 278 347 283 355
rect 285 347 290 368
rect 292 366 301 368
rect 292 364 297 366
rect 299 364 301 366
rect 292 358 301 364
rect 327 361 332 368
rect 325 359 332 361
rect 292 347 303 358
rect 257 343 260 345
rect 262 343 264 345
rect 257 341 264 343
rect 295 340 303 347
rect 305 356 312 358
rect 305 354 308 356
rect 310 354 312 356
rect 325 357 327 359
rect 329 357 332 359
rect 325 355 332 357
rect 305 349 312 354
rect 327 350 332 355
rect 334 366 342 368
rect 334 364 337 366
rect 339 364 342 366
rect 334 352 342 364
rect 344 352 349 368
rect 351 356 359 368
rect 351 354 354 356
rect 356 354 359 356
rect 351 352 359 354
rect 361 352 366 368
rect 368 366 375 368
rect 368 364 371 366
rect 373 364 375 366
rect 368 356 375 364
rect 401 361 406 368
rect 399 359 406 361
rect 399 357 401 359
rect 403 357 406 359
rect 368 352 374 356
rect 399 355 406 357
rect 334 350 339 352
rect 305 347 308 349
rect 310 347 312 349
rect 305 345 312 347
rect 305 340 310 345
rect 370 348 374 352
rect 401 350 406 355
rect 408 366 416 368
rect 408 364 411 366
rect 413 364 416 366
rect 408 352 416 364
rect 418 352 423 368
rect 425 356 433 368
rect 425 354 428 356
rect 430 354 433 356
rect 425 352 433 354
rect 435 352 440 368
rect 442 366 449 368
rect 442 364 445 366
rect 447 364 449 366
rect 442 356 449 364
rect 475 361 480 368
rect 473 359 480 361
rect 473 357 475 359
rect 477 357 480 359
rect 442 352 448 356
rect 473 355 480 357
rect 408 350 413 352
rect 370 340 376 348
rect 378 346 383 348
rect 378 344 385 346
rect 378 342 381 344
rect 383 342 385 344
rect 378 340 385 342
rect 444 348 448 352
rect 475 350 480 355
rect 482 366 490 368
rect 482 364 485 366
rect 487 364 490 366
rect 482 352 490 364
rect 492 352 497 368
rect 499 356 507 368
rect 499 354 502 356
rect 504 354 507 356
rect 499 352 507 354
rect 509 352 514 368
rect 516 366 523 368
rect 516 364 519 366
rect 521 364 523 366
rect 516 356 523 364
rect 516 352 522 356
rect 482 350 487 352
rect 444 340 450 348
rect 452 346 457 348
rect 452 344 459 346
rect 452 342 455 344
rect 457 342 459 344
rect 452 340 459 342
rect 518 348 522 352
rect 518 340 524 348
rect 526 346 531 348
rect 526 344 533 346
rect 526 342 529 344
rect 531 342 533 344
rect 526 340 533 342
rect -27 259 -22 264
rect -29 257 -22 259
rect -29 255 -27 257
rect -25 255 -22 257
rect -29 250 -22 255
rect -29 248 -27 250
rect -25 248 -22 250
rect -29 246 -22 248
rect -20 257 -12 264
rect 11 261 18 263
rect 11 259 13 261
rect 15 259 18 261
rect -20 246 -9 257
rect -18 240 -9 246
rect -18 238 -16 240
rect -14 238 -9 240
rect -18 236 -9 238
rect -7 236 -2 257
rect 0 249 5 257
rect 11 254 18 259
rect 11 252 13 254
rect 15 252 18 254
rect 11 250 18 252
rect 0 247 7 249
rect 0 245 3 247
rect 5 245 7 247
rect 13 245 18 250
rect 20 256 26 263
rect 59 261 66 263
rect 59 259 61 261
rect 63 259 66 261
rect 59 257 66 259
rect 20 249 28 256
rect 20 247 23 249
rect 25 247 28 249
rect 20 245 28 247
rect 0 243 7 245
rect 0 236 5 243
rect 22 243 28 245
rect 30 254 38 256
rect 30 252 33 254
rect 35 252 38 254
rect 30 247 38 252
rect 30 245 33 247
rect 35 245 38 247
rect 30 243 38 245
rect 40 247 47 256
rect 40 245 43 247
rect 45 245 47 247
rect 40 243 47 245
rect 61 236 66 257
rect 68 247 82 263
rect 68 245 71 247
rect 73 245 82 247
rect 84 261 92 263
rect 84 259 87 261
rect 89 259 92 261
rect 84 254 92 259
rect 84 252 87 254
rect 89 252 92 254
rect 84 245 92 252
rect 94 254 102 263
rect 94 252 97 254
rect 99 252 102 254
rect 94 245 102 252
rect 68 240 80 245
rect 68 238 71 240
rect 73 238 80 240
rect 68 236 80 238
rect 97 236 102 245
rect 104 248 109 263
rect 115 261 122 263
rect 115 259 117 261
rect 119 259 122 261
rect 115 254 122 259
rect 115 252 117 254
rect 119 252 122 254
rect 115 250 122 252
rect 104 246 111 248
rect 104 244 107 246
rect 109 244 111 246
rect 117 245 122 250
rect 124 256 130 263
rect 163 261 170 263
rect 163 259 165 261
rect 167 259 170 261
rect 163 257 170 259
rect 124 249 132 256
rect 124 247 127 249
rect 129 247 132 249
rect 124 245 132 247
rect 104 242 111 244
rect 104 236 109 242
rect 126 243 132 245
rect 134 254 142 256
rect 134 252 137 254
rect 139 252 142 254
rect 134 247 142 252
rect 134 245 137 247
rect 139 245 142 247
rect 134 243 142 245
rect 144 247 151 256
rect 144 245 147 247
rect 149 245 151 247
rect 144 243 151 245
rect 165 236 170 257
rect 172 247 186 263
rect 172 245 175 247
rect 177 245 186 247
rect 188 261 196 263
rect 188 259 191 261
rect 193 259 196 261
rect 188 254 196 259
rect 188 252 191 254
rect 193 252 196 254
rect 188 245 196 252
rect 198 254 206 263
rect 198 252 201 254
rect 203 252 206 254
rect 198 245 206 252
rect 172 240 184 245
rect 172 238 175 240
rect 177 238 184 240
rect 172 236 184 238
rect 201 236 206 245
rect 208 248 213 263
rect 249 256 255 263
rect 208 246 215 248
rect 208 244 211 246
rect 213 244 215 246
rect 208 242 215 244
rect 228 247 235 256
rect 228 245 230 247
rect 232 245 235 247
rect 228 243 235 245
rect 237 254 245 256
rect 237 252 240 254
rect 242 252 245 254
rect 237 247 245 252
rect 237 245 240 247
rect 242 245 245 247
rect 237 243 245 245
rect 247 249 255 256
rect 247 247 250 249
rect 252 247 255 249
rect 247 245 255 247
rect 257 261 264 263
rect 257 259 260 261
rect 262 259 264 261
rect 257 254 264 259
rect 295 257 303 264
rect 257 252 260 254
rect 262 252 264 254
rect 257 250 264 252
rect 257 245 262 250
rect 278 249 283 257
rect 276 247 283 249
rect 276 245 278 247
rect 280 245 283 247
rect 247 243 253 245
rect 208 236 213 242
rect 276 243 283 245
rect 278 236 283 243
rect 285 236 290 257
rect 292 246 303 257
rect 305 259 310 264
rect 305 257 312 259
rect 305 255 308 257
rect 310 255 312 257
rect 305 250 312 255
rect 305 248 308 250
rect 310 248 312 250
rect 327 249 332 254
rect 305 246 312 248
rect 325 247 332 249
rect 292 240 301 246
rect 325 245 327 247
rect 329 245 332 247
rect 325 243 332 245
rect 292 238 297 240
rect 299 238 301 240
rect 292 236 301 238
rect 327 236 332 243
rect 334 252 339 254
rect 370 256 376 264
rect 378 262 385 264
rect 378 260 381 262
rect 383 260 385 262
rect 378 258 385 260
rect 378 256 383 258
rect 370 252 374 256
rect 334 240 342 252
rect 334 238 337 240
rect 339 238 342 240
rect 334 236 342 238
rect 344 236 349 252
rect 351 250 359 252
rect 351 248 354 250
rect 356 248 359 250
rect 351 236 359 248
rect 361 236 366 252
rect 368 248 374 252
rect 401 249 406 254
rect 368 240 375 248
rect 399 247 406 249
rect 399 245 401 247
rect 403 245 406 247
rect 399 243 406 245
rect 368 238 371 240
rect 373 238 375 240
rect 368 236 375 238
rect 401 236 406 243
rect 408 252 413 254
rect 444 256 450 264
rect 452 262 459 264
rect 452 260 455 262
rect 457 260 459 262
rect 452 258 459 260
rect 452 256 457 258
rect 444 252 448 256
rect 408 240 416 252
rect 408 238 411 240
rect 413 238 416 240
rect 408 236 416 238
rect 418 236 423 252
rect 425 250 433 252
rect 425 248 428 250
rect 430 248 433 250
rect 425 236 433 248
rect 435 236 440 252
rect 442 248 448 252
rect 475 249 480 254
rect 442 240 449 248
rect 473 247 480 249
rect 473 245 475 247
rect 477 245 480 247
rect 473 243 480 245
rect 442 238 445 240
rect 447 238 449 240
rect 442 236 449 238
rect 475 236 480 243
rect 482 252 487 254
rect 518 256 524 264
rect 526 262 533 264
rect 526 260 529 262
rect 531 260 533 262
rect 526 258 533 260
rect 526 256 531 258
rect 518 252 522 256
rect 482 240 490 252
rect 482 238 485 240
rect 487 238 490 240
rect 482 236 490 238
rect 492 236 497 252
rect 499 250 507 252
rect 499 248 502 250
rect 504 248 507 250
rect 499 236 507 248
rect 509 236 514 252
rect 516 248 522 252
rect 516 240 523 248
rect 516 238 519 240
rect 521 238 523 240
rect 516 236 523 238
rect -18 222 -9 224
rect -18 220 -16 222
rect -14 220 -9 222
rect -18 214 -9 220
rect -29 212 -22 214
rect -29 210 -27 212
rect -25 210 -22 212
rect -29 205 -22 210
rect -29 203 -27 205
rect -25 203 -22 205
rect -29 201 -22 203
rect -27 196 -22 201
rect -20 203 -9 214
rect -7 203 -2 224
rect 0 217 5 224
rect 0 215 7 217
rect 22 215 28 217
rect 0 213 3 215
rect 5 213 7 215
rect 0 211 7 213
rect 0 203 5 211
rect 13 210 18 215
rect 11 208 18 210
rect 11 206 13 208
rect 15 206 18 208
rect -20 196 -12 203
rect 11 201 18 206
rect 11 199 13 201
rect 15 199 18 201
rect 11 197 18 199
rect 20 213 28 215
rect 20 211 23 213
rect 25 211 28 213
rect 20 204 28 211
rect 30 215 38 217
rect 30 213 33 215
rect 35 213 38 215
rect 30 208 38 213
rect 30 206 33 208
rect 35 206 38 208
rect 30 204 38 206
rect 40 215 47 217
rect 40 213 43 215
rect 45 213 47 215
rect 40 204 47 213
rect 20 197 26 204
rect 61 203 66 224
rect 59 201 66 203
rect 59 199 61 201
rect 63 199 66 201
rect 59 197 66 199
rect 68 222 80 224
rect 68 220 71 222
rect 73 220 80 222
rect 68 215 80 220
rect 97 215 102 224
rect 68 213 71 215
rect 73 213 82 215
rect 68 197 82 213
rect 84 208 92 215
rect 84 206 87 208
rect 89 206 92 208
rect 84 201 92 206
rect 84 199 87 201
rect 89 199 92 201
rect 84 197 92 199
rect 94 208 102 215
rect 94 206 97 208
rect 99 206 102 208
rect 94 197 102 206
rect 104 218 109 224
rect 104 216 111 218
rect 104 214 107 216
rect 109 214 111 216
rect 126 215 132 217
rect 104 212 111 214
rect 104 197 109 212
rect 117 210 122 215
rect 115 208 122 210
rect 115 206 117 208
rect 119 206 122 208
rect 115 201 122 206
rect 115 199 117 201
rect 119 199 122 201
rect 115 197 122 199
rect 124 213 132 215
rect 124 211 127 213
rect 129 211 132 213
rect 124 204 132 211
rect 134 215 142 217
rect 134 213 137 215
rect 139 213 142 215
rect 134 208 142 213
rect 134 206 137 208
rect 139 206 142 208
rect 134 204 142 206
rect 144 215 151 217
rect 144 213 147 215
rect 149 213 151 215
rect 144 204 151 213
rect 124 197 130 204
rect 165 203 170 224
rect 163 201 170 203
rect 163 199 165 201
rect 167 199 170 201
rect 163 197 170 199
rect 172 222 184 224
rect 172 220 175 222
rect 177 220 184 222
rect 172 215 184 220
rect 201 215 206 224
rect 172 213 175 215
rect 177 213 186 215
rect 172 197 186 213
rect 188 208 196 215
rect 188 206 191 208
rect 193 206 196 208
rect 188 201 196 206
rect 188 199 191 201
rect 193 199 196 201
rect 188 197 196 199
rect 198 208 206 215
rect 198 206 201 208
rect 203 206 206 208
rect 198 197 206 206
rect 208 218 213 224
rect 208 216 215 218
rect 208 214 211 216
rect 213 214 215 216
rect 208 212 215 214
rect 228 215 235 217
rect 228 213 230 215
rect 232 213 235 215
rect 208 197 213 212
rect 228 204 235 213
rect 237 215 245 217
rect 237 213 240 215
rect 242 213 245 215
rect 237 208 245 213
rect 237 206 240 208
rect 242 206 245 208
rect 237 204 245 206
rect 247 215 253 217
rect 278 217 283 224
rect 276 215 283 217
rect 247 213 255 215
rect 247 211 250 213
rect 252 211 255 213
rect 247 204 255 211
rect 249 197 255 204
rect 257 210 262 215
rect 276 213 278 215
rect 280 213 283 215
rect 276 211 283 213
rect 257 208 264 210
rect 257 206 260 208
rect 262 206 264 208
rect 257 201 264 206
rect 278 203 283 211
rect 285 203 290 224
rect 292 222 301 224
rect 292 220 297 222
rect 299 220 301 222
rect 292 214 301 220
rect 327 217 332 224
rect 325 215 332 217
rect 292 203 303 214
rect 257 199 260 201
rect 262 199 264 201
rect 257 197 264 199
rect 295 196 303 203
rect 305 212 312 214
rect 305 210 308 212
rect 310 210 312 212
rect 325 213 327 215
rect 329 213 332 215
rect 325 211 332 213
rect 305 205 312 210
rect 327 206 332 211
rect 334 222 342 224
rect 334 220 337 222
rect 339 220 342 222
rect 334 208 342 220
rect 344 208 349 224
rect 351 212 359 224
rect 351 210 354 212
rect 356 210 359 212
rect 351 208 359 210
rect 361 208 366 224
rect 368 222 375 224
rect 368 220 371 222
rect 373 220 375 222
rect 368 212 375 220
rect 401 217 406 224
rect 399 215 406 217
rect 399 213 401 215
rect 403 213 406 215
rect 368 208 374 212
rect 399 211 406 213
rect 334 206 339 208
rect 305 203 308 205
rect 310 203 312 205
rect 305 201 312 203
rect 305 196 310 201
rect 370 204 374 208
rect 401 206 406 211
rect 408 222 416 224
rect 408 220 411 222
rect 413 220 416 222
rect 408 208 416 220
rect 418 208 423 224
rect 425 212 433 224
rect 425 210 428 212
rect 430 210 433 212
rect 425 208 433 210
rect 435 208 440 224
rect 442 222 449 224
rect 442 220 445 222
rect 447 220 449 222
rect 442 212 449 220
rect 475 217 480 224
rect 473 215 480 217
rect 473 213 475 215
rect 477 213 480 215
rect 442 208 448 212
rect 473 211 480 213
rect 408 206 413 208
rect 370 196 376 204
rect 378 202 383 204
rect 378 200 385 202
rect 378 198 381 200
rect 383 198 385 200
rect 378 196 385 198
rect 444 204 448 208
rect 475 206 480 211
rect 482 222 490 224
rect 482 220 485 222
rect 487 220 490 222
rect 482 208 490 220
rect 492 208 497 224
rect 499 212 507 224
rect 499 210 502 212
rect 504 210 507 212
rect 499 208 507 210
rect 509 208 514 224
rect 516 222 523 224
rect 516 220 519 222
rect 521 220 523 222
rect 516 212 523 220
rect 516 208 522 212
rect 482 206 487 208
rect 444 196 450 204
rect 452 202 457 204
rect 452 200 459 202
rect 452 198 455 200
rect 457 198 459 200
rect 452 196 459 198
rect 518 204 522 208
rect 518 196 524 204
rect 526 202 531 204
rect 526 200 533 202
rect 526 198 529 200
rect 531 198 533 200
rect 526 196 533 198
<< alu1 >>
rect -33 441 537 446
rect -33 439 -26 441
rect -24 439 14 441
rect 16 439 24 441
rect 26 439 54 441
rect 56 439 107 441
rect 109 439 118 441
rect 120 439 128 441
rect 130 439 158 441
rect 160 439 211 441
rect 213 439 249 441
rect 251 439 259 441
rect 261 439 307 441
rect 309 439 537 441
rect -33 438 537 439
rect 11 429 23 433
rect 11 427 13 429
rect 15 427 23 429
rect 87 431 111 432
rect -29 424 -24 426
rect -29 422 -27 424
rect -25 422 -24 424
rect -29 420 -24 422
rect -29 401 -25 420
rect 3 416 7 425
rect -29 399 -27 401
rect -29 394 -25 399
rect -29 392 -27 394
rect -14 415 7 416
rect -14 413 -10 415
rect -8 413 4 415
rect 6 413 7 415
rect -14 412 7 413
rect -14 406 0 408
rect 2 406 7 408
rect -14 404 7 406
rect 3 402 7 404
rect 3 400 4 402
rect 6 400 7 402
rect 3 395 7 400
rect 11 407 15 427
rect 87 429 89 431
rect 91 429 111 431
rect 87 428 111 429
rect 35 424 40 425
rect 35 422 36 424
rect 38 422 40 424
rect 35 416 40 422
rect 11 405 16 407
rect 11 403 13 405
rect 15 403 16 405
rect 11 402 16 403
rect 11 400 12 402
rect 14 400 16 402
rect 11 398 16 400
rect 11 396 13 398
rect 15 396 16 398
rect 26 415 40 416
rect 26 413 30 415
rect 32 413 40 415
rect 26 412 40 413
rect 59 424 72 425
rect 59 422 61 424
rect 63 422 69 424
rect 71 422 72 424
rect 59 420 72 422
rect 59 419 69 420
rect 67 418 69 419
rect 71 418 72 420
rect 34 407 47 408
rect 34 405 40 407
rect 42 405 47 407
rect 34 404 47 405
rect 11 394 16 396
rect -29 388 -16 392
rect -29 387 -25 388
rect 43 400 47 404
rect 43 398 44 400
rect 46 398 47 400
rect 43 395 47 398
rect 51 407 56 409
rect 51 405 53 407
rect 55 405 56 407
rect 51 400 56 405
rect 67 411 72 418
rect 51 398 53 400
rect 55 398 56 400
rect 51 393 56 398
rect 51 387 63 393
rect 107 407 111 428
rect 107 405 108 407
rect 110 405 111 407
rect 107 400 111 405
rect 95 398 111 400
rect 95 396 97 398
rect 99 396 111 398
rect 95 395 111 396
rect 115 429 127 433
rect 115 427 117 429
rect 119 427 127 429
rect 191 431 215 432
rect 115 415 119 427
rect 191 429 193 431
rect 195 429 215 431
rect 191 428 215 429
rect 115 413 116 415
rect 118 413 119 415
rect 115 407 119 413
rect 139 424 144 425
rect 139 422 140 424
rect 142 422 144 424
rect 139 416 144 422
rect 115 405 120 407
rect 115 403 117 405
rect 119 403 120 405
rect 115 398 120 403
rect 115 396 117 398
rect 119 396 120 398
rect 130 415 144 416
rect 130 413 131 415
rect 133 413 134 415
rect 136 413 144 415
rect 130 412 144 413
rect 163 424 176 425
rect 163 422 165 424
rect 167 422 176 424
rect 163 420 176 422
rect 163 419 173 420
rect 171 418 173 419
rect 175 418 176 420
rect 138 407 151 408
rect 138 405 139 407
rect 141 405 144 407
rect 146 405 151 407
rect 138 404 151 405
rect 115 394 120 396
rect 147 400 151 404
rect 147 398 148 400
rect 150 398 151 400
rect 147 395 151 398
rect 155 407 160 409
rect 155 405 157 407
rect 159 405 160 407
rect 155 400 160 405
rect 171 411 176 418
rect 211 419 215 428
rect 211 417 212 419
rect 214 417 215 419
rect 155 398 157 400
rect 159 398 160 400
rect 155 393 160 398
rect 155 387 167 393
rect 211 400 215 417
rect 235 424 240 425
rect 235 422 237 424
rect 239 422 240 424
rect 235 416 240 422
rect 252 429 264 433
rect 252 427 260 429
rect 262 427 264 429
rect 235 415 249 416
rect 235 413 243 415
rect 245 413 249 415
rect 235 412 249 413
rect 199 398 215 400
rect 199 396 201 398
rect 203 396 215 398
rect 199 395 215 396
rect 228 407 241 408
rect 228 405 229 407
rect 231 405 233 407
rect 235 405 241 407
rect 228 404 241 405
rect 228 395 232 404
rect 260 410 264 427
rect 325 431 329 433
rect 325 429 330 431
rect 325 427 327 429
rect 329 427 330 429
rect 399 431 403 433
rect 276 424 280 425
rect 276 422 277 424
rect 279 422 280 424
rect 276 416 280 422
rect 276 415 297 416
rect 276 413 291 415
rect 293 413 297 415
rect 276 412 297 413
rect 307 424 312 426
rect 307 422 308 424
rect 310 422 312 424
rect 307 420 312 422
rect 260 408 261 410
rect 263 408 264 410
rect 260 407 264 408
rect 259 405 264 407
rect 259 403 260 405
rect 262 403 264 405
rect 259 398 264 403
rect 259 396 260 398
rect 262 396 264 398
rect 259 394 264 396
rect 276 407 281 408
rect 276 405 277 407
rect 279 406 281 407
rect 283 406 297 408
rect 279 405 297 406
rect 276 404 297 405
rect 276 395 280 404
rect 308 409 312 420
rect 308 407 309 409
rect 311 407 312 409
rect 308 401 312 407
rect 310 399 312 401
rect 308 394 312 399
rect 310 392 312 394
rect 299 388 312 392
rect 325 425 330 427
rect 325 417 329 425
rect 325 415 326 417
rect 328 415 329 417
rect 325 392 329 415
rect 334 409 336 411
rect 340 410 345 417
rect 340 408 341 410
rect 343 409 345 410
rect 343 408 353 409
rect 340 407 353 408
rect 340 405 341 407
rect 343 405 353 407
rect 340 403 353 405
rect 365 420 378 424
rect 365 418 368 420
rect 370 418 372 420
rect 365 417 372 418
rect 365 415 368 417
rect 370 415 372 417
rect 365 411 372 415
rect 370 404 372 406
rect 399 429 404 431
rect 399 427 401 429
rect 403 427 404 429
rect 473 431 477 433
rect 399 425 404 427
rect 399 413 403 425
rect 399 411 400 413
rect 402 411 403 413
rect 372 396 385 400
rect 380 395 385 396
rect 325 391 338 392
rect 380 393 381 395
rect 383 393 385 395
rect 325 389 327 391
rect 329 389 338 391
rect 325 388 338 389
rect 308 387 312 388
rect 380 387 385 393
rect 399 392 403 411
rect 415 415 421 417
rect 415 413 417 415
rect 419 413 421 415
rect 415 412 421 413
rect 408 409 410 411
rect 414 410 421 412
rect 414 408 415 410
rect 417 409 421 410
rect 417 408 427 409
rect 414 406 427 408
rect 415 403 427 406
rect 439 420 452 424
rect 439 415 445 420
rect 439 413 442 415
rect 444 413 445 415
rect 439 411 445 413
rect 444 404 446 406
rect 473 429 478 431
rect 473 427 475 429
rect 477 427 478 429
rect 473 425 478 427
rect 446 396 459 400
rect 454 395 459 396
rect 399 391 412 392
rect 454 393 455 395
rect 457 393 459 395
rect 399 389 401 391
rect 403 389 412 391
rect 399 388 412 389
rect 454 387 459 393
rect 473 392 477 425
rect 489 413 493 417
rect 482 409 484 411
rect 489 411 490 413
rect 492 411 493 413
rect 489 410 493 411
rect 491 409 493 410
rect 491 408 501 409
rect 489 403 501 408
rect 513 422 526 424
rect 513 420 516 422
rect 518 420 526 422
rect 513 415 519 420
rect 513 413 516 415
rect 518 413 519 415
rect 513 411 519 413
rect 518 404 520 406
rect 520 396 533 400
rect 528 395 533 396
rect 473 391 486 392
rect 528 393 529 395
rect 531 393 533 395
rect 473 389 475 391
rect 477 389 486 391
rect 473 388 486 389
rect 528 387 533 393
rect -33 381 537 382
rect -33 379 -26 381
rect -24 379 14 381
rect 16 379 87 381
rect 89 379 118 381
rect 120 379 191 381
rect 193 379 259 381
rect 261 379 307 381
rect 309 379 537 381
rect -33 369 537 379
rect -33 367 -26 369
rect -24 367 14 369
rect 16 367 87 369
rect 89 367 118 369
rect 120 367 191 369
rect 193 367 259 369
rect 261 367 307 369
rect 309 367 537 369
rect -33 366 537 367
rect -29 360 -25 361
rect -29 358 -28 360
rect -26 358 -16 360
rect -29 356 -16 358
rect -29 354 -27 356
rect -29 349 -25 354
rect -29 347 -27 349
rect -29 328 -25 347
rect 3 348 7 353
rect 3 346 4 348
rect 6 346 7 348
rect 3 344 7 346
rect -14 342 7 344
rect -14 340 0 342
rect 2 340 7 342
rect 11 352 16 354
rect 11 350 13 352
rect 15 350 16 352
rect 51 355 63 361
rect 11 348 16 350
rect 11 346 12 348
rect 14 346 16 348
rect 11 345 16 346
rect 11 343 13 345
rect 15 343 16 345
rect 11 341 16 343
rect 43 350 47 353
rect 43 348 44 350
rect 46 348 47 350
rect -29 326 -24 328
rect -29 324 -27 326
rect -25 324 -24 326
rect -29 322 -24 324
rect -14 335 7 336
rect -14 333 -10 335
rect -8 333 4 335
rect 6 333 7 335
rect -14 332 7 333
rect 3 323 7 332
rect 11 321 15 341
rect 43 344 47 348
rect 34 343 47 344
rect 34 341 40 343
rect 42 341 47 343
rect 34 340 47 341
rect 51 350 56 355
rect 51 348 53 350
rect 55 348 56 350
rect 51 343 56 348
rect 51 341 53 343
rect 55 341 56 343
rect 51 339 56 341
rect 26 335 40 336
rect 26 333 30 335
rect 32 333 40 335
rect 26 332 40 333
rect 11 319 13 321
rect 15 319 23 321
rect 11 315 23 319
rect 35 326 40 332
rect 35 324 36 326
rect 38 324 40 326
rect 35 323 40 324
rect 67 330 72 337
rect 95 352 111 353
rect 95 350 97 352
rect 99 350 111 352
rect 95 348 111 350
rect 107 343 111 348
rect 107 341 108 343
rect 110 341 111 343
rect 67 329 69 330
rect 59 328 69 329
rect 71 328 72 330
rect 59 326 72 328
rect 59 324 61 326
rect 63 324 72 326
rect 59 323 72 324
rect 107 320 111 341
rect 87 319 111 320
rect 87 317 89 319
rect 91 317 111 319
rect 87 316 111 317
rect 115 352 120 354
rect 115 350 117 352
rect 119 350 120 352
rect 155 355 167 361
rect 115 345 120 350
rect 115 343 117 345
rect 119 343 120 345
rect 115 341 120 343
rect 147 350 151 353
rect 147 348 148 350
rect 150 348 151 350
rect 115 335 119 341
rect 115 333 116 335
rect 118 333 119 335
rect 115 321 119 333
rect 147 344 151 348
rect 138 343 151 344
rect 138 341 139 343
rect 141 341 144 343
rect 146 341 151 343
rect 138 340 151 341
rect 155 350 160 355
rect 155 348 157 350
rect 159 348 160 350
rect 155 343 160 348
rect 155 341 157 343
rect 159 341 160 343
rect 155 339 160 341
rect 130 335 144 336
rect 130 333 131 335
rect 133 333 134 335
rect 136 333 144 335
rect 130 332 144 333
rect 115 319 117 321
rect 119 319 127 321
rect 115 315 127 319
rect 139 326 144 332
rect 139 324 140 326
rect 142 324 144 326
rect 139 323 144 324
rect 171 330 176 337
rect 199 352 215 353
rect 199 350 201 352
rect 203 350 215 352
rect 199 348 215 350
rect 171 329 173 330
rect 163 328 173 329
rect 175 328 176 330
rect 163 326 176 328
rect 163 324 165 326
rect 167 324 176 326
rect 163 323 176 324
rect 211 331 215 348
rect 228 344 232 353
rect 308 360 312 361
rect 299 356 312 360
rect 259 352 264 354
rect 228 343 241 344
rect 228 341 229 343
rect 231 341 233 343
rect 235 341 241 343
rect 228 340 241 341
rect 211 329 212 331
rect 214 329 215 331
rect 211 320 215 329
rect 235 335 249 336
rect 235 333 243 335
rect 245 333 249 335
rect 235 332 249 333
rect 259 350 260 352
rect 262 350 264 352
rect 259 345 264 350
rect 259 343 260 345
rect 262 343 264 345
rect 259 341 264 343
rect 235 326 240 332
rect 235 324 236 326
rect 238 324 240 326
rect 235 323 240 324
rect 260 340 264 341
rect 276 344 280 353
rect 276 343 297 344
rect 276 341 277 343
rect 279 342 297 343
rect 279 341 281 342
rect 276 340 281 341
rect 283 340 297 342
rect 260 338 261 340
rect 263 338 264 340
rect 260 321 264 338
rect 276 335 297 336
rect 276 333 291 335
rect 293 333 297 335
rect 276 332 297 333
rect 310 354 312 356
rect 308 349 312 354
rect 310 347 312 349
rect 276 326 280 332
rect 308 341 312 347
rect 308 339 309 341
rect 311 339 312 341
rect 308 328 312 339
rect 276 324 277 326
rect 279 324 280 326
rect 276 323 280 324
rect 307 326 312 328
rect 307 324 308 326
rect 310 324 312 326
rect 307 322 312 324
rect 325 359 338 360
rect 325 357 327 359
rect 329 357 338 359
rect 325 356 338 357
rect 325 333 329 356
rect 380 355 385 361
rect 380 353 381 355
rect 383 353 385 355
rect 325 331 326 333
rect 328 331 329 333
rect 380 352 385 353
rect 372 348 385 352
rect 399 359 412 360
rect 399 357 401 359
rect 403 357 412 359
rect 399 356 412 357
rect 334 337 336 339
rect 325 323 329 331
rect 340 343 353 345
rect 340 341 341 343
rect 343 341 353 343
rect 340 340 353 341
rect 340 338 341 340
rect 343 339 353 340
rect 370 342 372 344
rect 343 338 345 339
rect 340 331 345 338
rect 365 333 372 337
rect 365 331 368 333
rect 370 331 372 333
rect 365 330 372 331
rect 365 328 368 330
rect 370 328 372 330
rect 365 324 378 328
rect 191 319 215 320
rect 191 317 193 319
rect 195 317 215 319
rect 191 316 215 317
rect 252 319 260 321
rect 262 319 264 321
rect 252 315 264 319
rect 325 321 330 323
rect 325 319 327 321
rect 329 319 330 321
rect 325 317 330 319
rect 325 315 329 317
rect 399 337 403 356
rect 454 355 459 361
rect 454 353 455 355
rect 457 353 459 355
rect 399 335 400 337
rect 402 335 403 337
rect 399 323 403 335
rect 454 352 459 353
rect 446 348 459 352
rect 473 359 486 360
rect 473 357 475 359
rect 477 357 486 359
rect 473 356 486 357
rect 415 342 427 345
rect 408 337 410 339
rect 414 340 427 342
rect 414 338 415 340
rect 417 339 427 340
rect 444 342 446 344
rect 417 338 421 339
rect 414 336 421 338
rect 415 335 421 336
rect 415 333 417 335
rect 419 333 421 335
rect 415 331 421 333
rect 439 335 445 337
rect 439 333 442 335
rect 444 333 445 335
rect 439 328 445 333
rect 439 324 452 328
rect 399 321 404 323
rect 399 319 401 321
rect 403 319 404 321
rect 399 317 404 319
rect 399 315 403 317
rect 473 323 477 356
rect 528 355 533 361
rect 528 353 529 355
rect 531 353 533 355
rect 528 352 533 353
rect 520 348 533 352
rect 482 337 484 339
rect 489 340 501 345
rect 491 339 501 340
rect 518 342 520 344
rect 491 338 493 339
rect 489 337 493 338
rect 489 335 490 337
rect 492 335 493 337
rect 489 331 493 335
rect 513 335 519 337
rect 513 333 516 335
rect 518 333 519 335
rect 513 328 519 333
rect 513 326 516 328
rect 518 326 526 328
rect 513 324 526 326
rect 473 321 478 323
rect 473 319 475 321
rect 477 319 478 321
rect 473 317 478 319
rect 473 315 477 317
rect -33 309 537 310
rect -33 307 -26 309
rect -24 307 14 309
rect 16 307 24 309
rect 26 307 54 309
rect 56 307 107 309
rect 109 307 118 309
rect 120 307 128 309
rect 130 307 158 309
rect 160 307 211 309
rect 213 307 249 309
rect 251 307 259 309
rect 261 307 307 309
rect 309 307 537 309
rect -33 297 537 307
rect -33 295 -26 297
rect -24 295 14 297
rect 16 295 24 297
rect 26 295 54 297
rect 56 295 107 297
rect 109 295 118 297
rect 120 295 128 297
rect 130 295 158 297
rect 160 295 211 297
rect 213 295 249 297
rect 251 295 259 297
rect 261 295 307 297
rect 309 295 537 297
rect -33 294 537 295
rect 11 285 23 289
rect 11 283 13 285
rect 15 283 23 285
rect 87 287 111 288
rect -29 280 -24 282
rect -29 278 -27 280
rect -25 278 -24 280
rect -29 276 -24 278
rect -37 275 -25 276
rect -37 273 -36 275
rect -34 273 -25 275
rect -37 272 -25 273
rect -29 257 -25 272
rect 3 272 7 281
rect -29 255 -27 257
rect -29 250 -25 255
rect -29 248 -27 250
rect -14 271 7 272
rect -14 269 -10 271
rect -8 269 4 271
rect 6 269 7 271
rect -14 268 7 269
rect -14 262 0 264
rect 2 262 7 264
rect -14 260 7 262
rect 3 258 7 260
rect 3 256 4 258
rect 6 256 7 258
rect 3 251 7 256
rect 11 263 15 283
rect 87 285 89 287
rect 91 285 111 287
rect 87 284 111 285
rect 35 280 40 281
rect 35 278 36 280
rect 38 278 40 280
rect 35 272 40 278
rect 11 261 16 263
rect 11 259 13 261
rect 15 259 16 261
rect 11 258 16 259
rect 11 256 12 258
rect 14 256 16 258
rect 11 254 16 256
rect 11 252 13 254
rect 15 252 16 254
rect 26 271 40 272
rect 26 269 30 271
rect 32 269 40 271
rect 26 268 40 269
rect 59 280 72 281
rect 59 278 61 280
rect 63 278 69 280
rect 71 278 72 280
rect 59 276 72 278
rect 59 275 69 276
rect 67 274 69 275
rect 71 274 72 276
rect 34 263 47 264
rect 34 261 40 263
rect 42 261 47 263
rect 34 260 47 261
rect 11 250 16 252
rect -29 244 -16 248
rect -29 243 -25 244
rect 43 256 47 260
rect 43 254 44 256
rect 46 254 47 256
rect 43 251 47 254
rect 51 263 56 265
rect 51 261 53 263
rect 55 261 56 263
rect 51 256 56 261
rect 67 267 72 274
rect 51 254 53 256
rect 55 254 56 256
rect 51 249 56 254
rect 51 243 63 249
rect 107 263 111 284
rect 107 261 108 263
rect 110 261 111 263
rect 107 256 111 261
rect 95 254 111 256
rect 95 252 97 254
rect 99 252 111 254
rect 95 251 111 252
rect 115 285 127 289
rect 115 283 117 285
rect 119 283 127 285
rect 191 287 215 288
rect 115 271 119 283
rect 191 285 193 287
rect 195 285 215 287
rect 191 284 215 285
rect 115 269 116 271
rect 118 269 119 271
rect 115 263 119 269
rect 139 280 144 281
rect 139 278 140 280
rect 142 278 144 280
rect 139 272 144 278
rect 115 261 120 263
rect 115 259 117 261
rect 119 259 120 261
rect 115 254 120 259
rect 115 252 117 254
rect 119 252 120 254
rect 130 271 144 272
rect 130 269 131 271
rect 133 269 134 271
rect 136 269 144 271
rect 130 268 144 269
rect 163 280 176 281
rect 163 278 165 280
rect 167 278 176 280
rect 163 276 176 278
rect 163 275 173 276
rect 171 274 173 275
rect 175 274 176 276
rect 138 263 151 264
rect 138 261 139 263
rect 141 261 144 263
rect 146 261 151 263
rect 138 260 151 261
rect 115 250 120 252
rect 147 256 151 260
rect 147 254 148 256
rect 150 254 151 256
rect 147 251 151 254
rect 155 263 160 265
rect 155 261 157 263
rect 159 261 160 263
rect 155 256 160 261
rect 171 267 176 274
rect 211 275 215 284
rect 211 273 212 275
rect 214 273 215 275
rect 155 254 157 256
rect 159 254 160 256
rect 155 249 160 254
rect 155 243 167 249
rect 211 256 215 273
rect 235 280 240 281
rect 235 278 237 280
rect 239 278 240 280
rect 235 272 240 278
rect 252 285 264 289
rect 252 283 260 285
rect 262 283 264 285
rect 235 271 249 272
rect 235 269 243 271
rect 245 269 249 271
rect 235 268 249 269
rect 199 254 215 256
rect 199 252 201 254
rect 203 252 215 254
rect 199 251 215 252
rect 228 263 241 264
rect 228 261 229 263
rect 231 261 233 263
rect 235 261 241 263
rect 228 260 241 261
rect 228 251 232 260
rect 260 266 264 283
rect 325 287 329 289
rect 325 285 330 287
rect 325 283 327 285
rect 329 283 330 285
rect 399 287 403 289
rect 276 280 280 281
rect 276 278 277 280
rect 279 278 280 280
rect 276 272 280 278
rect 276 271 297 272
rect 276 269 291 271
rect 293 269 297 271
rect 276 268 297 269
rect 307 280 312 282
rect 307 278 308 280
rect 310 278 312 280
rect 307 276 312 278
rect 260 264 261 266
rect 263 264 264 266
rect 260 263 264 264
rect 259 261 264 263
rect 259 259 260 261
rect 262 259 264 261
rect 259 254 264 259
rect 259 252 260 254
rect 262 252 264 254
rect 259 250 264 252
rect 276 263 281 264
rect 276 261 277 263
rect 279 262 281 263
rect 283 262 297 264
rect 279 261 297 262
rect 276 260 297 261
rect 276 251 280 260
rect 308 265 312 276
rect 308 263 309 265
rect 311 263 312 265
rect 308 257 312 263
rect 310 255 312 257
rect 308 250 312 255
rect 310 248 312 250
rect 299 244 312 248
rect 325 281 330 283
rect 325 273 329 281
rect 325 271 326 273
rect 328 271 329 273
rect 325 248 329 271
rect 334 265 336 267
rect 340 266 345 273
rect 340 264 341 266
rect 343 265 345 266
rect 343 264 353 265
rect 340 263 353 264
rect 340 261 341 263
rect 343 261 353 263
rect 340 259 353 261
rect 365 276 378 280
rect 365 274 368 276
rect 370 274 372 276
rect 365 273 372 274
rect 365 271 368 273
rect 370 271 372 273
rect 365 267 372 271
rect 370 260 372 262
rect 399 285 404 287
rect 399 283 401 285
rect 403 283 404 285
rect 473 287 477 289
rect 399 281 404 283
rect 399 269 403 281
rect 399 267 400 269
rect 402 267 403 269
rect 372 252 385 256
rect 380 251 385 252
rect 325 247 338 248
rect 380 249 381 251
rect 383 249 385 251
rect 325 245 327 247
rect 329 245 338 247
rect 325 244 338 245
rect 308 243 312 244
rect 380 243 385 249
rect 399 248 403 267
rect 415 271 421 273
rect 415 269 417 271
rect 419 269 421 271
rect 415 268 421 269
rect 408 265 410 267
rect 414 266 421 268
rect 414 264 415 266
rect 417 265 421 266
rect 417 264 427 265
rect 414 262 427 264
rect 415 259 427 262
rect 439 276 452 280
rect 439 271 445 276
rect 439 269 442 271
rect 444 269 445 271
rect 439 267 445 269
rect 444 260 446 262
rect 473 285 478 287
rect 473 283 475 285
rect 477 283 478 285
rect 473 281 478 283
rect 446 252 459 256
rect 454 251 459 252
rect 399 247 412 248
rect 454 249 455 251
rect 457 249 459 251
rect 399 245 401 247
rect 403 245 412 247
rect 399 244 412 245
rect 454 243 459 249
rect 473 248 477 281
rect 489 269 493 273
rect 482 265 484 267
rect 489 267 490 269
rect 492 267 493 269
rect 489 266 493 267
rect 491 265 493 266
rect 491 264 501 265
rect 489 259 501 264
rect 513 278 526 280
rect 513 276 516 278
rect 518 276 526 278
rect 513 271 519 276
rect 513 269 516 271
rect 518 269 519 271
rect 513 267 519 269
rect 518 260 520 262
rect 520 252 533 256
rect 528 251 533 252
rect 473 247 486 248
rect 528 249 529 251
rect 531 249 533 251
rect 473 245 475 247
rect 477 245 486 247
rect 473 244 486 245
rect 528 243 533 249
rect -33 237 537 238
rect -33 235 -26 237
rect -24 235 14 237
rect 16 235 87 237
rect 89 235 118 237
rect 120 235 191 237
rect 193 235 259 237
rect 261 235 307 237
rect 309 235 537 237
rect -33 225 537 235
rect -33 223 -26 225
rect -24 223 14 225
rect 16 223 87 225
rect 89 223 118 225
rect 120 223 191 225
rect 193 223 259 225
rect 261 223 307 225
rect 309 223 537 225
rect -33 222 537 223
rect -29 216 -25 217
rect -29 214 -28 216
rect -26 214 -16 216
rect -29 212 -16 214
rect -29 210 -27 212
rect -29 205 -25 210
rect -29 203 -27 205
rect -29 184 -25 203
rect 3 204 7 209
rect 3 202 4 204
rect 6 202 7 204
rect 3 200 7 202
rect -14 198 7 200
rect -14 196 0 198
rect 2 196 7 198
rect 11 208 16 210
rect 11 206 13 208
rect 15 206 16 208
rect 51 211 63 217
rect 11 204 16 206
rect 11 202 12 204
rect 14 202 16 204
rect 11 201 16 202
rect 11 199 13 201
rect 15 199 16 201
rect 11 197 16 199
rect 43 206 47 209
rect 43 204 44 206
rect 46 204 47 206
rect -29 182 -24 184
rect -29 180 -27 182
rect -25 180 -24 182
rect -29 178 -24 180
rect -14 191 7 192
rect -14 189 -10 191
rect -8 189 4 191
rect 6 189 7 191
rect -14 188 7 189
rect 3 179 7 188
rect 11 177 15 197
rect 43 200 47 204
rect 34 199 47 200
rect 34 197 40 199
rect 42 197 47 199
rect 34 196 47 197
rect 51 206 56 211
rect 51 204 53 206
rect 55 204 56 206
rect 51 199 56 204
rect 51 197 53 199
rect 55 197 56 199
rect 51 195 56 197
rect 26 191 40 192
rect 26 189 30 191
rect 32 189 40 191
rect 26 188 40 189
rect 11 175 13 177
rect 15 175 23 177
rect 11 171 23 175
rect 35 182 40 188
rect 35 180 36 182
rect 38 180 40 182
rect 35 179 40 180
rect 67 186 72 193
rect 95 208 111 209
rect 95 206 97 208
rect 99 206 111 208
rect 95 204 111 206
rect 107 199 111 204
rect 107 197 108 199
rect 110 197 111 199
rect 67 185 69 186
rect 59 184 69 185
rect 71 184 72 186
rect 59 182 72 184
rect 59 180 61 182
rect 63 180 72 182
rect 59 179 72 180
rect 107 176 111 197
rect 87 175 111 176
rect 87 173 89 175
rect 91 173 111 175
rect 87 172 111 173
rect 115 208 120 210
rect 115 206 117 208
rect 119 206 120 208
rect 155 211 167 217
rect 115 201 120 206
rect 115 199 117 201
rect 119 199 120 201
rect 115 197 120 199
rect 147 206 151 209
rect 147 204 148 206
rect 150 204 151 206
rect 115 191 119 197
rect 115 189 116 191
rect 118 189 119 191
rect 115 177 119 189
rect 147 200 151 204
rect 138 199 151 200
rect 138 197 139 199
rect 141 197 144 199
rect 146 197 151 199
rect 138 196 151 197
rect 155 206 160 211
rect 155 204 157 206
rect 159 204 160 206
rect 155 199 160 204
rect 155 197 157 199
rect 159 197 160 199
rect 155 195 160 197
rect 130 191 144 192
rect 130 189 134 191
rect 136 189 144 191
rect 130 188 144 189
rect 115 175 117 177
rect 119 175 127 177
rect 115 171 127 175
rect 139 182 144 188
rect 139 180 140 182
rect 142 180 144 182
rect 139 179 144 180
rect 171 186 176 193
rect 199 208 215 209
rect 199 206 201 208
rect 203 206 215 208
rect 199 204 215 206
rect 171 185 173 186
rect 163 184 173 185
rect 175 184 176 186
rect 163 182 176 184
rect 163 180 165 182
rect 167 180 176 182
rect 163 179 176 180
rect 211 187 215 204
rect 228 200 232 209
rect 308 216 312 217
rect 299 212 312 216
rect 259 208 264 210
rect 228 199 241 200
rect 228 197 229 199
rect 231 197 233 199
rect 235 197 241 199
rect 228 196 241 197
rect 211 185 212 187
rect 214 185 215 187
rect 211 176 215 185
rect 235 191 249 192
rect 235 189 243 191
rect 245 189 249 191
rect 235 188 249 189
rect 259 206 260 208
rect 262 206 264 208
rect 259 201 264 206
rect 259 199 260 201
rect 262 199 264 201
rect 259 197 264 199
rect 235 182 240 188
rect 235 180 236 182
rect 238 180 240 182
rect 235 179 240 180
rect 260 196 264 197
rect 276 200 280 209
rect 276 199 297 200
rect 276 197 277 199
rect 279 198 297 199
rect 279 197 281 198
rect 276 196 281 197
rect 283 196 297 198
rect 260 194 261 196
rect 263 194 264 196
rect 260 177 264 194
rect 276 191 297 192
rect 276 189 291 191
rect 293 189 297 191
rect 276 188 297 189
rect 310 210 312 212
rect 308 205 312 210
rect 310 203 312 205
rect 276 182 280 188
rect 308 197 312 203
rect 308 195 309 197
rect 311 195 312 197
rect 308 184 312 195
rect 276 180 277 182
rect 279 180 280 182
rect 276 179 280 180
rect 307 182 312 184
rect 307 180 308 182
rect 310 180 312 182
rect 307 178 312 180
rect 325 215 338 216
rect 325 213 327 215
rect 329 213 338 215
rect 325 212 338 213
rect 325 189 329 212
rect 380 211 385 217
rect 380 209 381 211
rect 383 209 385 211
rect 325 187 326 189
rect 328 187 329 189
rect 380 208 385 209
rect 372 204 385 208
rect 399 215 412 216
rect 399 213 401 215
rect 403 213 412 215
rect 399 212 412 213
rect 334 193 336 195
rect 325 179 329 187
rect 340 199 353 201
rect 340 197 341 199
rect 343 197 353 199
rect 340 196 353 197
rect 340 194 341 196
rect 343 195 353 196
rect 370 198 372 200
rect 343 194 345 195
rect 340 187 345 194
rect 365 189 372 193
rect 365 187 368 189
rect 370 187 372 189
rect 365 186 372 187
rect 365 184 368 186
rect 370 184 372 186
rect 365 180 378 184
rect 191 175 215 176
rect 191 173 193 175
rect 195 173 215 175
rect 191 172 215 173
rect 252 175 260 177
rect 262 175 264 177
rect 252 171 264 175
rect 325 177 330 179
rect 325 175 327 177
rect 329 175 330 177
rect 325 173 330 175
rect 325 171 329 173
rect 399 193 403 212
rect 454 211 459 217
rect 454 209 455 211
rect 457 209 459 211
rect 399 191 400 193
rect 402 191 403 193
rect 399 179 403 191
rect 454 208 459 209
rect 446 204 459 208
rect 473 215 486 216
rect 473 213 475 215
rect 477 213 486 215
rect 473 212 486 213
rect 415 198 427 201
rect 408 193 410 195
rect 414 196 427 198
rect 414 194 415 196
rect 417 195 427 196
rect 444 198 446 200
rect 417 194 421 195
rect 414 192 421 194
rect 415 191 421 192
rect 415 189 417 191
rect 419 189 421 191
rect 415 187 421 189
rect 439 191 445 193
rect 439 189 442 191
rect 444 189 445 191
rect 439 184 445 189
rect 439 180 452 184
rect 399 177 404 179
rect 399 175 401 177
rect 403 175 404 177
rect 399 173 404 175
rect 399 171 403 173
rect 473 179 477 212
rect 528 211 533 217
rect 528 209 529 211
rect 531 209 533 211
rect 528 208 533 209
rect 520 204 533 208
rect 482 193 484 195
rect 489 196 501 201
rect 491 195 501 196
rect 518 198 520 200
rect 491 194 493 195
rect 489 193 493 194
rect 489 191 490 193
rect 492 191 493 193
rect 489 187 493 191
rect 513 191 519 193
rect 513 189 516 191
rect 518 189 519 191
rect 513 184 519 189
rect 513 182 516 184
rect 518 182 526 184
rect 513 180 526 182
rect 473 177 478 179
rect 473 175 475 177
rect 477 175 478 177
rect 473 173 478 175
rect 473 171 477 173
rect -33 165 537 166
rect -33 163 -26 165
rect -24 163 14 165
rect 16 163 24 165
rect 26 163 54 165
rect 56 163 107 165
rect 109 163 118 165
rect 120 163 128 165
rect 130 163 158 165
rect 160 163 211 165
rect 213 163 249 165
rect 251 163 259 165
rect 261 163 307 165
rect 309 163 537 165
rect -33 158 537 163
<< alu2 >>
rect 321 440 493 444
rect 35 424 72 425
rect 35 422 36 424
rect 38 422 61 424
rect 63 422 69 424
rect 71 422 72 424
rect 35 421 72 422
rect 139 424 171 425
rect 139 422 140 424
rect 142 422 165 424
rect 167 422 171 424
rect 35 420 67 421
rect 139 420 171 422
rect 236 424 240 425
rect 236 422 237 424
rect 239 422 240 424
rect 236 421 240 422
rect 276 424 280 425
rect 276 422 277 424
rect 279 422 280 424
rect 276 421 280 422
rect 211 419 224 420
rect 211 417 212 419
rect 214 417 224 419
rect 211 416 224 417
rect 3 415 119 416
rect 3 413 4 415
rect 6 413 116 415
rect 118 413 119 415
rect 3 412 119 413
rect 130 415 134 416
rect 130 413 131 415
rect 133 413 134 415
rect 130 412 134 413
rect 107 407 142 408
rect 107 405 108 407
rect 110 405 139 407
rect 141 405 142 407
rect 107 404 142 405
rect 3 402 16 403
rect 3 400 4 402
rect 6 400 12 402
rect 14 400 16 402
rect 3 398 16 400
rect 43 400 56 401
rect 43 398 44 400
rect 46 398 53 400
rect 55 398 56 400
rect 43 397 56 398
rect 147 400 160 401
rect 147 398 148 400
rect 150 398 157 400
rect 159 398 160 400
rect 147 397 160 398
rect 220 387 224 416
rect 321 418 325 440
rect 383 429 420 433
rect 321 417 329 418
rect 321 415 326 417
rect 328 415 329 417
rect 321 414 329 415
rect 367 417 371 420
rect 367 415 368 417
rect 370 415 371 417
rect 260 410 269 411
rect 340 410 344 411
rect 260 408 261 410
rect 263 408 269 410
rect 308 409 345 410
rect 228 407 232 408
rect 260 407 269 408
rect 228 405 229 407
rect 231 405 232 407
rect 228 404 232 405
rect 264 399 269 407
rect 276 407 280 408
rect 276 405 277 407
rect 279 405 280 407
rect 308 407 309 409
rect 311 407 345 409
rect 308 406 341 407
rect 276 404 280 405
rect 340 405 341 406
rect 343 405 345 407
rect 340 403 345 405
rect 367 399 371 415
rect 264 395 371 399
rect 383 387 387 429
rect 416 415 420 429
rect 220 383 387 387
rect 393 413 403 414
rect 393 411 400 413
rect 402 411 403 413
rect 393 410 403 411
rect 416 413 417 415
rect 419 413 420 415
rect 393 380 397 410
rect 416 407 420 413
rect 489 413 493 440
rect 489 411 490 413
rect 492 411 493 413
rect 489 406 493 411
rect 515 422 519 423
rect 515 420 516 422
rect 518 420 519 422
rect 515 380 519 420
rect 393 376 519 380
rect 393 368 519 372
rect 220 361 387 365
rect -29 360 -25 361
rect -29 358 -28 360
rect -26 358 -25 360
rect -29 357 -25 358
rect 43 350 56 351
rect 3 348 16 350
rect 3 346 4 348
rect 6 346 12 348
rect 14 346 16 348
rect 43 348 44 350
rect 46 348 53 350
rect 55 348 56 350
rect 43 347 56 348
rect 147 350 160 351
rect 147 348 148 350
rect 150 348 157 350
rect 159 348 160 350
rect 147 347 160 348
rect 3 345 16 346
rect 107 343 142 344
rect 107 341 108 343
rect 110 341 139 343
rect 141 341 142 343
rect 107 340 142 341
rect 3 335 119 336
rect 3 333 4 335
rect 6 333 116 335
rect 118 333 119 335
rect 3 332 119 333
rect 130 335 134 336
rect 130 333 131 335
rect 133 333 134 335
rect 130 332 134 333
rect 220 332 224 361
rect 264 349 371 353
rect 228 343 232 344
rect 228 341 229 343
rect 231 341 232 343
rect 264 341 269 349
rect 228 340 232 341
rect 260 340 269 341
rect 276 343 280 344
rect 276 341 277 343
rect 279 341 280 343
rect 340 343 345 345
rect 340 342 341 343
rect 276 340 280 341
rect 308 341 341 342
rect 343 341 345 343
rect 260 338 261 340
rect 263 338 269 340
rect 308 339 309 341
rect 311 339 345 341
rect 308 338 345 339
rect 260 337 269 338
rect 340 337 344 338
rect 211 331 224 332
rect 211 329 212 331
rect 214 329 224 331
rect 211 328 224 329
rect 321 333 329 334
rect 321 331 326 333
rect 328 331 329 333
rect 321 330 329 331
rect 367 333 371 349
rect 367 331 368 333
rect 370 331 371 333
rect 35 326 67 328
rect 35 324 36 326
rect 38 324 61 326
rect 63 324 67 326
rect 35 323 67 324
rect 139 326 171 328
rect 139 324 140 326
rect 142 324 165 326
rect 167 324 171 326
rect 139 323 171 324
rect 235 326 239 327
rect 235 324 236 326
rect 238 324 239 326
rect 235 323 239 324
rect 276 326 280 327
rect 276 324 277 326
rect 279 324 280 326
rect 276 323 280 324
rect 321 308 325 330
rect 367 328 371 331
rect 383 319 387 361
rect 393 338 397 368
rect 393 337 403 338
rect 393 335 400 337
rect 402 335 403 337
rect 393 334 403 335
rect 416 335 420 341
rect 416 333 417 335
rect 419 333 420 335
rect 416 319 420 333
rect 383 315 420 319
rect 489 337 493 342
rect 489 335 490 337
rect 492 335 493 337
rect 489 308 493 335
rect 515 328 519 368
rect 515 326 516 328
rect 518 326 519 328
rect 515 325 519 326
rect 321 304 493 308
rect 321 296 493 300
rect 35 280 72 281
rect 35 278 36 280
rect 38 278 61 280
rect 63 278 69 280
rect 71 278 72 280
rect 35 277 72 278
rect 139 280 171 281
rect 139 278 140 280
rect 142 278 165 280
rect 167 278 171 280
rect 35 276 67 277
rect 139 276 171 278
rect 236 280 240 281
rect 236 278 237 280
rect 239 278 240 280
rect 236 277 240 278
rect 276 280 280 281
rect 276 278 277 280
rect 279 278 280 280
rect 276 277 280 278
rect -37 275 -33 276
rect -37 273 -36 275
rect -34 273 -33 275
rect -37 272 -33 273
rect 211 275 224 276
rect 211 273 212 275
rect 214 273 224 275
rect 211 272 224 273
rect 3 271 119 272
rect 3 269 4 271
rect 6 269 116 271
rect 118 269 119 271
rect 3 268 119 269
rect 130 271 134 272
rect 130 269 131 271
rect 133 269 134 271
rect 130 268 134 269
rect 107 263 142 264
rect 107 261 108 263
rect 110 261 139 263
rect 141 261 142 263
rect 107 260 142 261
rect 3 258 16 259
rect 3 256 4 258
rect 6 256 12 258
rect 14 256 16 258
rect 3 254 16 256
rect 43 256 56 257
rect 43 254 44 256
rect 46 254 53 256
rect 55 254 56 256
rect 43 253 56 254
rect 147 256 160 257
rect 147 254 148 256
rect 150 254 157 256
rect 159 254 160 256
rect 147 253 160 254
rect 220 243 224 272
rect 321 274 325 296
rect 383 285 420 289
rect 321 273 329 274
rect 321 271 326 273
rect 328 271 329 273
rect 321 270 329 271
rect 367 273 371 276
rect 367 271 368 273
rect 370 271 371 273
rect 260 266 269 267
rect 340 266 344 267
rect 260 264 261 266
rect 263 264 269 266
rect 308 265 345 266
rect 228 263 232 264
rect 260 263 269 264
rect 228 261 229 263
rect 231 261 232 263
rect 228 260 232 261
rect 264 255 269 263
rect 276 263 280 264
rect 276 261 277 263
rect 279 261 280 263
rect 308 263 309 265
rect 311 263 345 265
rect 308 262 341 263
rect 276 260 280 261
rect 340 261 341 262
rect 343 261 345 263
rect 340 259 345 261
rect 367 255 371 271
rect 264 251 371 255
rect 383 243 387 285
rect 416 271 420 285
rect 220 239 387 243
rect 393 269 403 270
rect 393 267 400 269
rect 402 267 403 269
rect 393 266 403 267
rect 416 269 417 271
rect 419 269 420 271
rect 393 236 397 266
rect 416 263 420 269
rect 489 269 493 296
rect 489 267 490 269
rect 492 267 493 269
rect 489 262 493 267
rect 515 278 519 279
rect 515 276 516 278
rect 518 276 519 278
rect 515 236 519 276
rect 393 232 519 236
rect 393 224 519 228
rect 220 217 387 221
rect -29 216 -25 217
rect -29 214 -28 216
rect -26 214 -25 216
rect -29 213 -25 214
rect 43 206 56 207
rect 3 204 16 206
rect 3 202 4 204
rect 6 202 12 204
rect 14 202 16 204
rect 43 204 44 206
rect 46 204 53 206
rect 55 204 56 206
rect 43 203 56 204
rect 147 206 160 207
rect 147 204 148 206
rect 150 204 157 206
rect 159 204 160 206
rect 147 203 160 204
rect 3 201 16 202
rect 107 199 142 200
rect 107 197 108 199
rect 110 197 139 199
rect 141 197 142 199
rect 107 196 142 197
rect 3 191 119 192
rect 3 189 4 191
rect 6 189 116 191
rect 118 189 119 191
rect 3 188 119 189
rect 220 188 224 217
rect 264 205 371 209
rect 228 199 232 200
rect 228 197 229 199
rect 231 197 232 199
rect 264 197 269 205
rect 228 196 232 197
rect 260 196 269 197
rect 276 199 280 200
rect 276 197 277 199
rect 279 197 280 199
rect 340 199 345 201
rect 340 198 341 199
rect 276 196 280 197
rect 308 197 341 198
rect 343 197 345 199
rect 260 194 261 196
rect 263 194 269 196
rect 308 195 309 197
rect 311 195 345 197
rect 308 194 345 195
rect 260 193 269 194
rect 340 193 344 194
rect 211 187 224 188
rect 211 185 212 187
rect 214 185 224 187
rect 211 184 224 185
rect 321 189 329 190
rect 321 187 326 189
rect 328 187 329 189
rect 321 186 329 187
rect 367 189 371 205
rect 367 187 368 189
rect 370 187 371 189
rect 35 182 67 184
rect 35 180 36 182
rect 38 180 61 182
rect 63 180 67 182
rect 35 179 67 180
rect 139 182 171 184
rect 139 180 140 182
rect 142 180 165 182
rect 167 180 171 182
rect 139 179 171 180
rect 235 182 239 183
rect 235 180 236 182
rect 238 180 239 182
rect 235 179 239 180
rect 276 182 280 183
rect 276 180 277 182
rect 279 180 280 182
rect 276 179 280 180
rect 321 164 325 186
rect 367 184 371 187
rect 383 175 387 217
rect 393 194 397 224
rect 393 193 403 194
rect 393 191 400 193
rect 402 191 403 193
rect 393 190 403 191
rect 416 191 420 197
rect 416 189 417 191
rect 419 189 420 191
rect 416 175 420 189
rect 383 171 420 175
rect 489 193 493 198
rect 489 191 490 193
rect 492 191 493 193
rect 489 164 493 191
rect 515 184 519 224
rect 515 182 516 184
rect 518 182 519 184
rect 515 181 519 182
rect 321 160 493 164
<< alu3 >>
rect 67 424 280 425
rect 67 422 69 424
rect 71 422 237 424
rect 239 422 277 424
rect 279 422 280 424
rect 67 421 280 422
rect -29 415 136 416
rect -29 413 131 415
rect 133 413 136 415
rect -29 412 136 413
rect -29 360 -25 412
rect 51 407 280 408
rect 51 405 229 407
rect 231 405 277 407
rect 279 405 280 407
rect 51 404 280 405
rect 51 400 56 404
rect 51 398 53 400
rect 55 398 56 400
rect 51 397 56 398
rect -29 358 -28 360
rect -26 358 -25 360
rect -29 354 -25 358
rect 51 350 232 351
rect 51 348 53 350
rect 55 348 232 350
rect 51 347 232 348
rect 228 344 232 347
rect 228 343 280 344
rect 228 341 229 343
rect 231 341 277 343
rect 279 341 280 343
rect 228 340 280 341
rect 132 336 136 337
rect -29 335 136 336
rect -29 333 131 335
rect 133 333 136 335
rect -29 332 136 333
rect -29 305 -25 332
rect 60 326 280 327
rect 60 324 61 326
rect 63 324 236 326
rect 238 324 277 326
rect 279 324 280 326
rect 60 323 280 324
rect -37 301 -25 305
rect -37 275 -33 301
rect 67 280 280 281
rect 67 278 69 280
rect 71 278 237 280
rect 239 278 277 280
rect 279 278 280 280
rect 67 277 280 278
rect -37 273 -36 275
rect -34 273 -33 275
rect -37 272 -33 273
rect -29 271 136 272
rect -29 269 131 271
rect 133 269 136 271
rect -29 268 136 269
rect -29 216 -25 268
rect 51 263 280 264
rect 51 261 229 263
rect 231 261 277 263
rect 279 261 280 263
rect 51 260 280 261
rect 51 256 56 260
rect 51 254 53 256
rect 55 254 56 256
rect 51 253 56 254
rect -29 214 -28 216
rect -26 214 -25 216
rect -29 210 -25 214
rect 51 206 232 207
rect 51 204 53 206
rect 55 204 232 206
rect 51 203 232 204
rect 228 200 232 203
rect 228 199 280 200
rect 228 197 229 199
rect 231 197 277 199
rect 279 197 280 199
rect 228 196 280 197
rect 60 182 280 183
rect 60 180 61 182
rect 63 180 236 182
rect 238 180 277 182
rect 279 180 280 182
rect 60 179 280 180
<< ptie >>
rect -28 441 -22 443
rect -28 439 -26 441
rect -24 439 -22 441
rect 12 441 18 443
rect 12 439 14 441
rect 16 439 18 441
rect -28 437 -22 439
rect 12 437 18 439
rect 52 441 58 443
rect 52 439 54 441
rect 56 439 58 441
rect 52 437 58 439
rect 116 441 122 443
rect 116 439 118 441
rect 120 439 122 441
rect 116 437 122 439
rect 156 441 162 443
rect 156 439 158 441
rect 160 439 162 441
rect 156 437 162 439
rect 257 441 263 443
rect 257 439 259 441
rect 261 439 263 441
rect 305 441 311 443
rect 305 439 307 441
rect 309 439 311 441
rect 257 437 263 439
rect 305 437 311 439
rect -28 309 -22 311
rect 12 309 18 311
rect -28 307 -26 309
rect -24 307 -22 309
rect -28 305 -22 307
rect 12 307 14 309
rect 16 307 18 309
rect 12 305 18 307
rect 52 309 58 311
rect 52 307 54 309
rect 56 307 58 309
rect 52 305 58 307
rect 116 309 122 311
rect 116 307 118 309
rect 120 307 122 309
rect 116 305 122 307
rect 156 309 162 311
rect 156 307 158 309
rect 160 307 162 309
rect 156 305 162 307
rect 257 309 263 311
rect 305 309 311 311
rect 257 307 259 309
rect 261 307 263 309
rect 257 305 263 307
rect 305 307 307 309
rect 309 307 311 309
rect 305 305 311 307
rect -28 297 -22 299
rect -28 295 -26 297
rect -24 295 -22 297
rect 12 297 18 299
rect 12 295 14 297
rect 16 295 18 297
rect -28 293 -22 295
rect 12 293 18 295
rect 52 297 58 299
rect 52 295 54 297
rect 56 295 58 297
rect 52 293 58 295
rect 116 297 122 299
rect 116 295 118 297
rect 120 295 122 297
rect 116 293 122 295
rect 156 297 162 299
rect 156 295 158 297
rect 160 295 162 297
rect 156 293 162 295
rect 257 297 263 299
rect 257 295 259 297
rect 261 295 263 297
rect 305 297 311 299
rect 305 295 307 297
rect 309 295 311 297
rect 257 293 263 295
rect 305 293 311 295
rect -28 165 -22 167
rect 12 165 18 167
rect -28 163 -26 165
rect -24 163 -22 165
rect -28 161 -22 163
rect 12 163 14 165
rect 16 163 18 165
rect 12 161 18 163
rect 52 165 58 167
rect 52 163 54 165
rect 56 163 58 165
rect 52 161 58 163
rect 116 165 122 167
rect 116 163 118 165
rect 120 163 122 165
rect 116 161 122 163
rect 156 165 162 167
rect 156 163 158 165
rect 160 163 162 165
rect 156 161 162 163
rect 257 165 263 167
rect 305 165 311 167
rect 257 163 259 165
rect 261 163 263 165
rect 257 161 263 163
rect 305 163 307 165
rect 309 163 311 165
rect 305 161 311 163
<< ntie >>
rect -28 381 -22 383
rect -28 379 -26 381
rect -24 379 -22 381
rect 12 381 18 383
rect -28 377 -22 379
rect 12 379 14 381
rect 16 379 18 381
rect 85 381 91 383
rect 12 377 18 379
rect 85 379 87 381
rect 89 379 91 381
rect 116 381 122 383
rect 85 377 91 379
rect 116 379 118 381
rect 120 379 122 381
rect 189 381 195 383
rect 116 377 122 379
rect 189 379 191 381
rect 193 379 195 381
rect 257 381 263 383
rect 189 377 195 379
rect 257 379 259 381
rect 261 379 263 381
rect 305 381 311 383
rect 257 377 263 379
rect 305 379 307 381
rect 309 379 311 381
rect 305 377 311 379
rect -28 369 -22 371
rect -28 367 -26 369
rect -24 367 -22 369
rect 12 369 18 371
rect -28 365 -22 367
rect 12 367 14 369
rect 16 367 18 369
rect 85 369 91 371
rect 12 365 18 367
rect 85 367 87 369
rect 89 367 91 369
rect 116 369 122 371
rect 85 365 91 367
rect 116 367 118 369
rect 120 367 122 369
rect 189 369 195 371
rect 116 365 122 367
rect 189 367 191 369
rect 193 367 195 369
rect 257 369 263 371
rect 189 365 195 367
rect 257 367 259 369
rect 261 367 263 369
rect 305 369 311 371
rect 257 365 263 367
rect 305 367 307 369
rect 309 367 311 369
rect 305 365 311 367
rect -28 237 -22 239
rect -28 235 -26 237
rect -24 235 -22 237
rect 12 237 18 239
rect -28 233 -22 235
rect 12 235 14 237
rect 16 235 18 237
rect 85 237 91 239
rect 12 233 18 235
rect 85 235 87 237
rect 89 235 91 237
rect 116 237 122 239
rect 85 233 91 235
rect 116 235 118 237
rect 120 235 122 237
rect 189 237 195 239
rect 116 233 122 235
rect 189 235 191 237
rect 193 235 195 237
rect 257 237 263 239
rect 189 233 195 235
rect 257 235 259 237
rect 261 235 263 237
rect 305 237 311 239
rect 257 233 263 235
rect 305 235 307 237
rect 309 235 311 237
rect 305 233 311 235
rect -28 225 -22 227
rect -28 223 -26 225
rect -24 223 -22 225
rect 12 225 18 227
rect -28 221 -22 223
rect 12 223 14 225
rect 16 223 18 225
rect 85 225 91 227
rect 12 221 18 223
rect 85 223 87 225
rect 89 223 91 225
rect 116 225 122 227
rect 85 221 91 223
rect 116 223 118 225
rect 120 223 122 225
rect 189 225 195 227
rect 116 221 122 223
rect 189 223 191 225
rect 193 223 195 225
rect 257 225 263 227
rect 189 221 195 223
rect 257 223 259 225
rect 261 223 263 225
rect 305 225 311 227
rect 257 221 263 223
rect 305 223 307 225
rect 309 223 311 225
rect 305 221 311 223
<< nmos >>
rect -22 420 -20 429
rect -12 420 -10 426
rect -2 420 0 426
rect 18 422 20 431
rect 31 422 33 433
rect 38 422 40 433
rect 58 420 60 429
rect 74 425 76 434
rect 84 425 86 434
rect 94 425 96 437
rect 101 425 103 437
rect 122 422 124 431
rect 135 422 137 433
rect 142 422 144 433
rect 162 420 164 429
rect 178 425 180 434
rect 188 425 190 434
rect 198 425 200 437
rect 205 425 207 437
rect 235 422 237 433
rect 242 422 244 433
rect 255 422 257 431
rect 283 420 285 426
rect 293 420 295 426
rect 303 420 305 429
rect 332 425 334 434
rect 342 426 344 434
rect 349 426 351 434
rect 359 426 361 434
rect 366 426 368 434
rect 376 426 378 432
rect 406 425 408 434
rect 416 426 418 434
rect 423 426 425 434
rect 433 426 435 434
rect 440 426 442 434
rect 450 426 452 432
rect 480 425 482 434
rect 490 426 492 434
rect 497 426 499 434
rect 507 426 509 434
rect 514 426 516 434
rect 524 426 526 432
rect -22 319 -20 328
rect -12 322 -10 328
rect -2 322 0 328
rect 18 317 20 326
rect 31 315 33 326
rect 38 315 40 326
rect 58 319 60 328
rect 74 314 76 323
rect 84 314 86 323
rect 94 311 96 323
rect 101 311 103 323
rect 122 317 124 326
rect 135 315 137 326
rect 142 315 144 326
rect 162 319 164 328
rect 178 314 180 323
rect 188 314 190 323
rect 198 311 200 323
rect 205 311 207 323
rect 235 315 237 326
rect 242 315 244 326
rect 255 317 257 326
rect 283 322 285 328
rect 293 322 295 328
rect 303 319 305 328
rect 332 314 334 323
rect 342 314 344 322
rect 349 314 351 322
rect 359 314 361 322
rect 366 314 368 322
rect 376 316 378 322
rect 406 314 408 323
rect 416 314 418 322
rect 423 314 425 322
rect 433 314 435 322
rect 440 314 442 322
rect 450 316 452 322
rect 480 314 482 323
rect 490 314 492 322
rect 497 314 499 322
rect 507 314 509 322
rect 514 314 516 322
rect 524 316 526 322
rect -22 276 -20 285
rect -12 276 -10 282
rect -2 276 0 282
rect 18 278 20 287
rect 31 278 33 289
rect 38 278 40 289
rect 58 276 60 285
rect 74 281 76 290
rect 84 281 86 290
rect 94 281 96 293
rect 101 281 103 293
rect 122 278 124 287
rect 135 278 137 289
rect 142 278 144 289
rect 162 276 164 285
rect 178 281 180 290
rect 188 281 190 290
rect 198 281 200 293
rect 205 281 207 293
rect 235 278 237 289
rect 242 278 244 289
rect 255 278 257 287
rect 283 276 285 282
rect 293 276 295 282
rect 303 276 305 285
rect 332 281 334 290
rect 342 282 344 290
rect 349 282 351 290
rect 359 282 361 290
rect 366 282 368 290
rect 376 282 378 288
rect 406 281 408 290
rect 416 282 418 290
rect 423 282 425 290
rect 433 282 435 290
rect 440 282 442 290
rect 450 282 452 288
rect 480 281 482 290
rect 490 282 492 290
rect 497 282 499 290
rect 507 282 509 290
rect 514 282 516 290
rect 524 282 526 288
rect -22 175 -20 184
rect -12 178 -10 184
rect -2 178 0 184
rect 18 173 20 182
rect 31 171 33 182
rect 38 171 40 182
rect 58 175 60 184
rect 74 170 76 179
rect 84 170 86 179
rect 94 167 96 179
rect 101 167 103 179
rect 122 173 124 182
rect 135 171 137 182
rect 142 171 144 182
rect 162 175 164 184
rect 178 170 180 179
rect 188 170 190 179
rect 198 167 200 179
rect 205 167 207 179
rect 235 171 237 182
rect 242 171 244 182
rect 255 173 257 182
rect 283 178 285 184
rect 293 178 295 184
rect 303 175 305 184
rect 332 170 334 179
rect 342 170 344 178
rect 349 170 351 178
rect 359 170 361 178
rect 366 170 368 178
rect 376 172 378 178
rect 406 170 408 179
rect 416 170 418 178
rect 423 170 425 178
rect 433 170 435 178
rect 440 170 442 178
rect 450 172 452 178
rect 480 170 482 179
rect 490 170 492 178
rect 497 170 499 178
rect 507 170 509 178
rect 514 170 516 178
rect 524 172 526 178
<< pmos >>
rect -22 390 -20 408
rect -9 380 -7 401
rect -2 380 0 401
rect 18 389 20 407
rect 28 387 30 400
rect 38 387 40 400
rect 66 380 68 407
rect 82 389 84 407
rect 92 389 94 407
rect 102 380 104 407
rect 122 389 124 407
rect 132 387 134 400
rect 142 387 144 400
rect 170 380 172 407
rect 186 389 188 407
rect 196 389 198 407
rect 206 380 208 407
rect 235 387 237 400
rect 245 387 247 400
rect 255 389 257 407
rect 283 380 285 401
rect 290 380 292 401
rect 303 390 305 408
rect 332 380 334 398
rect 376 400 378 408
rect 342 380 344 396
rect 349 380 351 396
rect 359 380 361 396
rect 366 380 368 396
rect 406 380 408 398
rect 450 400 452 408
rect 416 380 418 396
rect 423 380 425 396
rect 433 380 435 396
rect 440 380 442 396
rect 480 380 482 398
rect 524 400 526 408
rect 490 380 492 396
rect 497 380 499 396
rect 507 380 509 396
rect 514 380 516 396
rect -22 340 -20 358
rect -9 347 -7 368
rect -2 347 0 368
rect 18 341 20 359
rect 28 348 30 361
rect 38 348 40 361
rect 66 341 68 368
rect 82 341 84 359
rect 92 341 94 359
rect 102 341 104 368
rect 122 341 124 359
rect 132 348 134 361
rect 142 348 144 361
rect 170 341 172 368
rect 186 341 188 359
rect 196 341 198 359
rect 206 341 208 368
rect 235 348 237 361
rect 245 348 247 361
rect 255 341 257 359
rect 283 347 285 368
rect 290 347 292 368
rect 303 340 305 358
rect 332 350 334 368
rect 342 352 344 368
rect 349 352 351 368
rect 359 352 361 368
rect 366 352 368 368
rect 406 350 408 368
rect 416 352 418 368
rect 423 352 425 368
rect 433 352 435 368
rect 440 352 442 368
rect 376 340 378 348
rect 480 350 482 368
rect 490 352 492 368
rect 497 352 499 368
rect 507 352 509 368
rect 514 352 516 368
rect 450 340 452 348
rect 524 340 526 348
rect -22 246 -20 264
rect -9 236 -7 257
rect -2 236 0 257
rect 18 245 20 263
rect 28 243 30 256
rect 38 243 40 256
rect 66 236 68 263
rect 82 245 84 263
rect 92 245 94 263
rect 102 236 104 263
rect 122 245 124 263
rect 132 243 134 256
rect 142 243 144 256
rect 170 236 172 263
rect 186 245 188 263
rect 196 245 198 263
rect 206 236 208 263
rect 235 243 237 256
rect 245 243 247 256
rect 255 245 257 263
rect 283 236 285 257
rect 290 236 292 257
rect 303 246 305 264
rect 332 236 334 254
rect 376 256 378 264
rect 342 236 344 252
rect 349 236 351 252
rect 359 236 361 252
rect 366 236 368 252
rect 406 236 408 254
rect 450 256 452 264
rect 416 236 418 252
rect 423 236 425 252
rect 433 236 435 252
rect 440 236 442 252
rect 480 236 482 254
rect 524 256 526 264
rect 490 236 492 252
rect 497 236 499 252
rect 507 236 509 252
rect 514 236 516 252
rect -22 196 -20 214
rect -9 203 -7 224
rect -2 203 0 224
rect 18 197 20 215
rect 28 204 30 217
rect 38 204 40 217
rect 66 197 68 224
rect 82 197 84 215
rect 92 197 94 215
rect 102 197 104 224
rect 122 197 124 215
rect 132 204 134 217
rect 142 204 144 217
rect 170 197 172 224
rect 186 197 188 215
rect 196 197 198 215
rect 206 197 208 224
rect 235 204 237 217
rect 245 204 247 217
rect 255 197 257 215
rect 283 203 285 224
rect 290 203 292 224
rect 303 196 305 214
rect 332 206 334 224
rect 342 208 344 224
rect 349 208 351 224
rect 359 208 361 224
rect 366 208 368 224
rect 406 206 408 224
rect 416 208 418 224
rect 423 208 425 224
rect 433 208 435 224
rect 440 208 442 224
rect 376 196 378 204
rect 480 206 482 224
rect 490 208 492 224
rect 497 208 499 224
rect 507 208 509 224
rect 514 208 516 224
rect 450 196 452 204
rect 524 196 526 204
<< polyct0 >>
rect -20 413 -18 415
rect 20 413 22 415
rect 90 413 92 415
rect 100 412 102 414
rect 124 413 126 415
rect 194 413 196 415
rect 204 412 206 414
rect 253 413 255 415
rect 333 418 335 420
rect 301 413 303 415
rect 351 419 353 421
rect 358 403 360 405
rect 407 418 409 420
rect 425 419 427 421
rect 432 403 434 405
rect 481 418 483 420
rect 499 419 501 421
rect 506 403 508 405
rect -20 333 -18 335
rect 20 333 22 335
rect 90 333 92 335
rect 100 334 102 336
rect 124 333 126 335
rect 194 333 196 335
rect 204 334 206 336
rect 253 333 255 335
rect 301 333 303 335
rect 358 343 360 345
rect 333 328 335 330
rect 351 327 353 329
rect 432 343 434 345
rect 407 328 409 330
rect 425 327 427 329
rect 506 343 508 345
rect 481 328 483 330
rect 499 327 501 329
rect -20 269 -18 271
rect 20 269 22 271
rect 90 269 92 271
rect 100 268 102 270
rect 124 269 126 271
rect 194 269 196 271
rect 204 268 206 270
rect 253 269 255 271
rect 333 274 335 276
rect 301 269 303 271
rect 351 275 353 277
rect 358 259 360 261
rect 407 274 409 276
rect 425 275 427 277
rect 432 259 434 261
rect 481 274 483 276
rect 499 275 501 277
rect 506 259 508 261
rect -20 189 -18 191
rect 20 189 22 191
rect 90 189 92 191
rect 100 190 102 192
rect 124 189 126 191
rect 194 189 196 191
rect 204 190 206 192
rect 253 189 255 191
rect 301 189 303 191
rect 358 199 360 201
rect 333 184 335 186
rect 351 183 353 185
rect 432 199 434 201
rect 407 184 409 186
rect 425 183 427 185
rect 506 199 508 201
rect 481 184 483 186
rect 499 183 501 185
<< polyct1 >>
rect -10 413 -8 415
rect 30 413 32 415
rect 0 406 2 408
rect 69 418 71 420
rect 40 405 42 407
rect 134 413 136 415
rect 53 405 55 407
rect 173 418 175 420
rect 144 405 146 407
rect 243 413 245 415
rect 157 405 159 407
rect 233 405 235 407
rect 291 413 293 415
rect 281 406 283 408
rect 341 408 343 410
rect 368 418 370 420
rect 415 408 417 410
rect 442 413 444 415
rect 381 393 383 395
rect 489 408 491 410
rect 516 413 518 415
rect 455 393 457 395
rect 529 393 531 395
rect 0 340 2 342
rect -10 333 -8 335
rect 40 341 42 343
rect 53 341 55 343
rect 30 333 32 335
rect 144 341 146 343
rect 157 341 159 343
rect 233 341 235 343
rect 69 328 71 330
rect 134 333 136 335
rect 173 328 175 330
rect 281 340 283 342
rect 243 333 245 335
rect 381 353 383 355
rect 291 333 293 335
rect 341 338 343 340
rect 455 353 457 355
rect 368 328 370 330
rect 415 338 417 340
rect 529 353 531 355
rect 442 333 444 335
rect 489 338 491 340
rect 516 333 518 335
rect -10 269 -8 271
rect 30 269 32 271
rect 0 262 2 264
rect 69 274 71 276
rect 40 261 42 263
rect 134 269 136 271
rect 53 261 55 263
rect 173 274 175 276
rect 144 261 146 263
rect 243 269 245 271
rect 157 261 159 263
rect 233 261 235 263
rect 291 269 293 271
rect 281 262 283 264
rect 341 264 343 266
rect 368 274 370 276
rect 415 264 417 266
rect 442 269 444 271
rect 381 249 383 251
rect 489 264 491 266
rect 516 269 518 271
rect 455 249 457 251
rect 529 249 531 251
rect 0 196 2 198
rect -10 189 -8 191
rect 40 197 42 199
rect 53 197 55 199
rect 30 189 32 191
rect 144 197 146 199
rect 157 197 159 199
rect 233 197 235 199
rect 69 184 71 186
rect 134 189 136 191
rect 173 184 175 186
rect 281 196 283 198
rect 243 189 245 191
rect 381 209 383 211
rect 291 189 293 191
rect 341 194 343 196
rect 455 209 457 211
rect 368 184 370 186
rect 415 194 417 196
rect 529 209 531 211
rect 442 189 444 191
rect 489 194 491 196
rect 516 189 518 191
<< ndifct0 >>
rect -16 435 -14 437
rect 3 435 5 437
rect -7 422 -5 424
rect 43 429 45 431
rect 67 430 69 432
rect 53 422 55 424
rect 79 427 81 429
rect 147 429 149 431
rect 171 430 173 432
rect 157 422 159 424
rect 183 427 185 429
rect 278 435 280 437
rect 230 429 232 431
rect 297 435 299 437
rect 288 422 290 424
rect 337 430 339 432
rect 354 430 356 432
rect 371 428 373 430
rect 381 428 383 430
rect 411 430 413 432
rect 428 430 430 432
rect 445 428 447 430
rect 455 428 457 430
rect 485 430 487 432
rect 502 430 504 432
rect 519 428 521 430
rect 529 428 531 430
rect -7 324 -5 326
rect -16 311 -14 313
rect 53 324 55 326
rect 43 317 45 319
rect 67 316 69 318
rect 3 311 5 313
rect 79 319 81 321
rect 157 324 159 326
rect 147 317 149 319
rect 171 316 173 318
rect 183 319 185 321
rect 230 317 232 319
rect 288 324 290 326
rect 278 311 280 313
rect 337 316 339 318
rect 354 316 356 318
rect 371 318 373 320
rect 381 318 383 320
rect 297 311 299 313
rect 411 316 413 318
rect 428 316 430 318
rect 445 318 447 320
rect 455 318 457 320
rect 485 316 487 318
rect 502 316 504 318
rect 519 318 521 320
rect 529 318 531 320
rect -16 291 -14 293
rect 3 291 5 293
rect -7 278 -5 280
rect 43 285 45 287
rect 67 286 69 288
rect 53 278 55 280
rect 79 283 81 285
rect 147 285 149 287
rect 171 286 173 288
rect 157 278 159 280
rect 183 283 185 285
rect 278 291 280 293
rect 230 285 232 287
rect 297 291 299 293
rect 288 278 290 280
rect 337 286 339 288
rect 354 286 356 288
rect 371 284 373 286
rect 381 284 383 286
rect 411 286 413 288
rect 428 286 430 288
rect 445 284 447 286
rect 455 284 457 286
rect 485 286 487 288
rect 502 286 504 288
rect 519 284 521 286
rect 529 284 531 286
rect -7 180 -5 182
rect -16 167 -14 169
rect 53 180 55 182
rect 43 173 45 175
rect 67 172 69 174
rect 3 167 5 169
rect 79 175 81 177
rect 157 180 159 182
rect 147 173 149 175
rect 171 172 173 174
rect 183 175 185 177
rect 230 173 232 175
rect 288 180 290 182
rect 278 167 280 169
rect 337 172 339 174
rect 354 172 356 174
rect 371 174 373 176
rect 381 174 383 176
rect 297 167 299 169
rect 411 172 413 174
rect 428 172 430 174
rect 445 174 447 176
rect 455 174 457 176
rect 485 172 487 174
rect 502 172 504 174
rect 519 174 521 176
rect 529 174 531 176
<< ndifct1 >>
rect 24 439 26 441
rect -27 422 -25 424
rect 107 439 109 441
rect 128 439 130 441
rect 13 427 15 429
rect 89 429 91 431
rect 211 439 213 441
rect 249 439 251 441
rect 117 427 119 429
rect 193 429 195 431
rect 260 427 262 429
rect 327 427 329 429
rect 401 427 403 429
rect 308 422 310 424
rect 475 427 477 429
rect -27 324 -25 326
rect 13 319 15 321
rect 89 317 91 319
rect 24 307 26 309
rect 117 319 119 321
rect 107 307 109 309
rect 193 317 195 319
rect 128 307 130 309
rect 260 319 262 321
rect 211 307 213 309
rect 308 324 310 326
rect 327 319 329 321
rect 249 307 251 309
rect 401 319 403 321
rect 475 319 477 321
rect 24 295 26 297
rect -27 278 -25 280
rect 107 295 109 297
rect 128 295 130 297
rect 13 283 15 285
rect 89 285 91 287
rect 211 295 213 297
rect 249 295 251 297
rect 117 283 119 285
rect 193 285 195 287
rect 260 283 262 285
rect 327 283 329 285
rect 401 283 403 285
rect 308 278 310 280
rect 475 283 477 285
rect -27 180 -25 182
rect 13 175 15 177
rect 89 173 91 175
rect 24 163 26 165
rect 117 175 119 177
rect 107 163 109 165
rect 193 173 195 175
rect 128 163 130 165
rect 260 175 262 177
rect 211 163 213 165
rect 308 180 310 182
rect 327 175 329 177
rect 249 163 251 165
rect 401 175 403 177
rect 475 175 477 177
<< ntiect1 >>
rect -26 379 -24 381
rect 14 379 16 381
rect 87 379 89 381
rect 118 379 120 381
rect 191 379 193 381
rect 259 379 261 381
rect 307 379 309 381
rect -26 367 -24 369
rect 14 367 16 369
rect 87 367 89 369
rect 118 367 120 369
rect 191 367 193 369
rect 259 367 261 369
rect 307 367 309 369
rect -26 235 -24 237
rect 14 235 16 237
rect 87 235 89 237
rect 118 235 120 237
rect 191 235 193 237
rect 259 235 261 237
rect 307 235 309 237
rect -26 223 -24 225
rect 14 223 16 225
rect 87 223 89 225
rect 118 223 120 225
rect 191 223 193 225
rect 259 223 261 225
rect 307 223 309 225
<< ptiect1 >>
rect -26 439 -24 441
rect 14 439 16 441
rect 54 439 56 441
rect 118 439 120 441
rect 158 439 160 441
rect 259 439 261 441
rect 307 439 309 441
rect -26 307 -24 309
rect 14 307 16 309
rect 54 307 56 309
rect 118 307 120 309
rect 158 307 160 309
rect 259 307 261 309
rect 307 307 309 309
rect -26 295 -24 297
rect 14 295 16 297
rect 54 295 56 297
rect 118 295 120 297
rect 158 295 160 297
rect 259 295 261 297
rect 307 295 309 297
rect -26 163 -24 165
rect 14 163 16 165
rect 54 163 56 165
rect 118 163 120 165
rect 158 163 160 165
rect 259 163 261 165
rect 307 163 309 165
<< pdifct0 >>
rect -16 382 -14 384
rect 3 389 5 391
rect 61 403 63 405
rect 23 391 25 393
rect 33 396 35 398
rect 33 389 35 391
rect 43 389 45 391
rect 71 389 73 391
rect 87 403 89 405
rect 87 396 89 398
rect 71 382 73 384
rect 107 388 109 390
rect 165 403 167 405
rect 127 391 129 393
rect 137 396 139 398
rect 137 389 139 391
rect 147 389 149 391
rect 175 389 177 391
rect 191 403 193 405
rect 191 396 193 398
rect 175 382 177 384
rect 211 388 213 390
rect 230 389 232 391
rect 240 396 242 398
rect 240 389 242 391
rect 250 391 252 393
rect 278 389 280 391
rect 297 382 299 384
rect 381 404 383 406
rect 337 382 339 384
rect 354 392 356 394
rect 371 382 373 384
rect 455 404 457 406
rect 411 382 413 384
rect 428 392 430 394
rect 445 382 447 384
rect 529 404 531 406
rect 485 382 487 384
rect 502 392 504 394
rect 519 382 521 384
rect -16 364 -14 366
rect 3 357 5 359
rect 23 355 25 357
rect 33 357 35 359
rect 33 350 35 352
rect 43 357 45 359
rect 61 343 63 345
rect 71 364 73 366
rect 71 357 73 359
rect 87 350 89 352
rect 87 343 89 345
rect 107 358 109 360
rect 127 355 129 357
rect 137 357 139 359
rect 137 350 139 352
rect 147 357 149 359
rect 165 343 167 345
rect 175 364 177 366
rect 175 357 177 359
rect 191 350 193 352
rect 191 343 193 345
rect 211 358 213 360
rect 230 357 232 359
rect 240 357 242 359
rect 240 350 242 352
rect 250 355 252 357
rect 278 357 280 359
rect 297 364 299 366
rect 337 364 339 366
rect 354 354 356 356
rect 371 364 373 366
rect 411 364 413 366
rect 428 354 430 356
rect 445 364 447 366
rect 381 342 383 344
rect 485 364 487 366
rect 502 354 504 356
rect 519 364 521 366
rect 455 342 457 344
rect 529 342 531 344
rect -16 238 -14 240
rect 3 245 5 247
rect 61 259 63 261
rect 23 247 25 249
rect 33 252 35 254
rect 33 245 35 247
rect 43 245 45 247
rect 71 245 73 247
rect 87 259 89 261
rect 87 252 89 254
rect 71 238 73 240
rect 107 244 109 246
rect 165 259 167 261
rect 127 247 129 249
rect 137 252 139 254
rect 137 245 139 247
rect 147 245 149 247
rect 175 245 177 247
rect 191 259 193 261
rect 191 252 193 254
rect 175 238 177 240
rect 211 244 213 246
rect 230 245 232 247
rect 240 252 242 254
rect 240 245 242 247
rect 250 247 252 249
rect 278 245 280 247
rect 297 238 299 240
rect 381 260 383 262
rect 337 238 339 240
rect 354 248 356 250
rect 371 238 373 240
rect 455 260 457 262
rect 411 238 413 240
rect 428 248 430 250
rect 445 238 447 240
rect 529 260 531 262
rect 485 238 487 240
rect 502 248 504 250
rect 519 238 521 240
rect -16 220 -14 222
rect 3 213 5 215
rect 23 211 25 213
rect 33 213 35 215
rect 33 206 35 208
rect 43 213 45 215
rect 61 199 63 201
rect 71 220 73 222
rect 71 213 73 215
rect 87 206 89 208
rect 87 199 89 201
rect 107 214 109 216
rect 127 211 129 213
rect 137 213 139 215
rect 137 206 139 208
rect 147 213 149 215
rect 165 199 167 201
rect 175 220 177 222
rect 175 213 177 215
rect 191 206 193 208
rect 191 199 193 201
rect 211 214 213 216
rect 230 213 232 215
rect 240 213 242 215
rect 240 206 242 208
rect 250 211 252 213
rect 278 213 280 215
rect 297 220 299 222
rect 337 220 339 222
rect 354 210 356 212
rect 371 220 373 222
rect 411 220 413 222
rect 428 210 430 212
rect 445 220 447 222
rect 381 198 383 200
rect 485 220 487 222
rect 502 210 504 212
rect 519 220 521 222
rect 455 198 457 200
rect 529 198 531 200
<< pdifct1 >>
rect -27 399 -25 401
rect -27 392 -25 394
rect 13 403 15 405
rect 13 396 15 398
rect 97 396 99 398
rect 117 403 119 405
rect 117 396 119 398
rect 201 396 203 398
rect 260 403 262 405
rect 260 396 262 398
rect 308 399 310 401
rect 308 392 310 394
rect 327 389 329 391
rect 401 389 403 391
rect 475 389 477 391
rect -27 354 -25 356
rect -27 347 -25 349
rect 13 350 15 352
rect 13 343 15 345
rect 97 350 99 352
rect 117 350 119 352
rect 117 343 119 345
rect 201 350 203 352
rect 260 350 262 352
rect 260 343 262 345
rect 308 354 310 356
rect 327 357 329 359
rect 401 357 403 359
rect 308 347 310 349
rect 475 357 477 359
rect -27 255 -25 257
rect -27 248 -25 250
rect 13 259 15 261
rect 13 252 15 254
rect 97 252 99 254
rect 117 259 119 261
rect 117 252 119 254
rect 201 252 203 254
rect 260 259 262 261
rect 260 252 262 254
rect 308 255 310 257
rect 308 248 310 250
rect 327 245 329 247
rect 401 245 403 247
rect 475 245 477 247
rect -27 210 -25 212
rect -27 203 -25 205
rect 13 206 15 208
rect 13 199 15 201
rect 97 206 99 208
rect 117 206 119 208
rect 117 199 119 201
rect 201 206 203 208
rect 260 206 262 208
rect 260 199 262 201
rect 308 210 310 212
rect 327 213 329 215
rect 401 213 403 215
rect 308 203 310 205
rect 475 213 477 215
<< alu0 >>
rect -18 437 -12 438
rect -18 435 -16 437
rect -14 435 -12 437
rect -18 434 -12 435
rect 1 437 7 438
rect 1 435 3 437
rect 5 435 7 437
rect 1 434 7 435
rect 65 432 71 438
rect 27 431 47 432
rect 27 429 43 431
rect 45 429 47 431
rect 65 430 67 432
rect 69 430 71 432
rect 65 429 71 430
rect 78 429 82 431
rect 27 428 47 429
rect -21 424 -3 425
rect -21 422 -7 424
rect -5 422 -3 424
rect -21 421 -3 422
rect -21 415 -17 421
rect -21 413 -20 415
rect -18 413 -17 415
rect -25 392 -24 403
rect -21 400 -17 413
rect -2 408 4 409
rect -21 396 -6 400
rect -10 392 -6 396
rect 15 425 16 427
rect 27 424 31 428
rect 78 427 79 429
rect 81 427 82 429
rect 19 420 31 424
rect 19 415 23 420
rect 19 413 20 415
rect 22 413 23 415
rect 19 401 23 413
rect 52 424 56 426
rect 52 422 53 424
rect 55 422 56 424
rect 52 416 56 422
rect 78 424 82 427
rect 78 420 102 424
rect 52 412 63 416
rect 19 398 36 401
rect 19 397 33 398
rect 32 396 33 397
rect 35 396 36 398
rect 21 393 27 394
rect -10 391 7 392
rect -10 389 3 391
rect 5 389 7 391
rect -10 388 7 389
rect 21 391 23 393
rect 25 391 27 393
rect -18 384 -12 385
rect -18 382 -16 384
rect -14 382 -12 384
rect 21 382 27 391
rect 32 391 36 396
rect 59 406 63 412
rect 98 416 102 420
rect 78 415 94 416
rect 78 413 90 415
rect 92 413 94 415
rect 78 412 94 413
rect 98 414 103 416
rect 98 412 100 414
rect 102 412 103 414
rect 78 406 82 412
rect 98 410 103 412
rect 98 408 102 410
rect 59 405 82 406
rect 59 403 61 405
rect 63 403 82 405
rect 59 402 82 403
rect 32 389 33 391
rect 35 389 36 391
rect 32 387 36 389
rect 41 391 47 392
rect 41 389 43 391
rect 45 389 47 391
rect 41 382 47 389
rect 70 391 74 393
rect 70 389 71 391
rect 73 389 74 391
rect 70 384 74 389
rect 78 391 82 402
rect 86 405 102 408
rect 86 403 87 405
rect 89 404 102 405
rect 89 403 90 404
rect 86 398 90 403
rect 86 396 87 398
rect 89 396 90 398
rect 86 394 90 396
rect 169 432 175 438
rect 276 437 282 438
rect 276 435 278 437
rect 280 435 282 437
rect 276 434 282 435
rect 295 437 301 438
rect 295 435 297 437
rect 299 435 301 437
rect 295 434 301 435
rect 131 431 151 432
rect 131 429 147 431
rect 149 429 151 431
rect 169 430 171 432
rect 173 430 175 432
rect 169 429 175 430
rect 182 429 186 431
rect 131 428 151 429
rect 119 425 120 427
rect 131 424 135 428
rect 182 427 183 429
rect 185 427 186 429
rect 228 431 248 432
rect 228 429 230 431
rect 232 429 248 431
rect 228 428 248 429
rect 123 420 135 424
rect 123 415 127 420
rect 123 413 124 415
rect 126 413 127 415
rect 123 401 127 413
rect 156 424 160 426
rect 156 422 157 424
rect 159 422 160 424
rect 156 416 160 422
rect 182 424 186 427
rect 182 420 206 424
rect 156 412 167 416
rect 123 398 140 401
rect 123 397 137 398
rect 136 396 137 397
rect 139 396 140 398
rect 125 393 131 394
rect 125 391 127 393
rect 129 391 131 393
rect 78 390 111 391
rect 78 388 107 390
rect 109 388 111 390
rect 78 387 111 388
rect 70 382 71 384
rect 73 382 74 384
rect 125 382 131 391
rect 136 391 140 396
rect 163 406 167 412
rect 202 416 206 420
rect 182 415 198 416
rect 182 413 194 415
rect 196 413 198 415
rect 182 412 198 413
rect 202 414 207 416
rect 202 412 204 414
rect 206 412 207 414
rect 182 406 186 412
rect 202 410 207 412
rect 202 408 206 410
rect 163 405 186 406
rect 163 403 165 405
rect 167 403 186 405
rect 163 402 186 403
rect 136 389 137 391
rect 139 389 140 391
rect 136 387 140 389
rect 145 391 151 392
rect 145 389 147 391
rect 149 389 151 391
rect 145 382 151 389
rect 174 391 178 393
rect 174 389 175 391
rect 177 389 178 391
rect 174 384 178 389
rect 182 391 186 402
rect 190 405 206 408
rect 190 403 191 405
rect 193 404 206 405
rect 193 403 194 404
rect 190 398 194 403
rect 244 424 248 428
rect 259 425 260 427
rect 244 420 256 424
rect 252 415 256 420
rect 252 413 253 415
rect 255 413 256 415
rect 190 396 191 398
rect 193 396 194 398
rect 190 394 194 396
rect 252 401 256 413
rect 336 432 340 438
rect 336 430 337 432
rect 339 430 340 432
rect 336 428 340 430
rect 343 432 358 433
rect 343 430 354 432
rect 356 430 358 432
rect 343 429 358 430
rect 369 430 375 438
rect 410 432 414 438
rect 286 424 304 425
rect 286 422 288 424
rect 290 422 304 424
rect 286 421 304 422
rect 300 415 304 421
rect 300 413 301 415
rect 303 413 304 415
rect 279 408 285 409
rect 239 398 256 401
rect 239 396 240 398
rect 242 397 256 398
rect 242 396 243 397
rect 228 391 234 392
rect 182 390 215 391
rect 182 388 211 390
rect 213 388 215 390
rect 182 387 215 388
rect 228 389 230 391
rect 232 389 234 391
rect 174 382 175 384
rect 177 382 178 384
rect 228 382 234 389
rect 239 391 243 396
rect 300 400 304 413
rect 289 396 304 400
rect 239 389 240 391
rect 242 389 243 391
rect 239 387 243 389
rect 248 393 254 394
rect 248 391 250 393
rect 252 391 254 393
rect 289 392 293 396
rect 307 392 308 403
rect 248 382 254 391
rect 276 391 293 392
rect 276 389 278 391
rect 280 389 293 391
rect 276 388 293 389
rect 343 424 347 429
rect 369 428 371 430
rect 373 428 375 430
rect 369 427 375 428
rect 379 430 385 431
rect 379 428 381 430
rect 383 428 385 430
rect 379 427 385 428
rect 333 422 347 424
rect 332 420 347 422
rect 350 421 361 423
rect 332 418 333 420
rect 335 418 337 420
rect 332 416 337 418
rect 350 419 351 421
rect 353 419 361 421
rect 350 417 361 419
rect 333 411 337 416
rect 333 409 334 411
rect 336 409 337 411
rect 333 399 337 409
rect 357 407 361 417
rect 381 407 385 427
rect 357 406 385 407
rect 357 405 370 406
rect 357 403 358 405
rect 360 404 370 405
rect 372 404 381 406
rect 383 404 385 406
rect 360 403 385 404
rect 410 430 411 432
rect 413 430 414 432
rect 410 428 414 430
rect 417 432 432 433
rect 417 430 428 432
rect 430 430 432 432
rect 417 429 432 430
rect 443 430 449 438
rect 484 432 488 438
rect 417 424 421 429
rect 443 428 445 430
rect 447 428 449 430
rect 443 427 449 428
rect 453 430 459 431
rect 453 428 455 430
rect 457 428 459 430
rect 453 427 459 428
rect 407 422 421 424
rect 406 420 421 422
rect 424 421 435 423
rect 406 418 407 420
rect 409 418 411 420
rect 406 416 411 418
rect 424 419 425 421
rect 427 419 435 421
rect 424 417 435 419
rect 357 401 361 403
rect 333 395 349 399
rect 345 394 358 395
rect 345 392 354 394
rect 356 392 358 394
rect 345 391 358 392
rect 407 411 411 416
rect 407 409 408 411
rect 410 409 411 411
rect 407 399 411 409
rect 431 407 435 417
rect 455 407 459 427
rect 431 406 459 407
rect 431 405 444 406
rect 431 403 432 405
rect 434 404 444 405
rect 446 404 455 406
rect 457 404 459 406
rect 434 403 459 404
rect 484 430 485 432
rect 487 430 488 432
rect 484 428 488 430
rect 491 432 506 433
rect 491 430 502 432
rect 504 430 506 432
rect 491 429 506 430
rect 517 430 523 438
rect 431 401 435 403
rect 407 395 423 399
rect 419 394 432 395
rect 419 392 428 394
rect 430 392 432 394
rect 419 391 432 392
rect 491 424 495 429
rect 517 428 519 430
rect 521 428 523 430
rect 517 427 523 428
rect 527 430 533 431
rect 527 428 529 430
rect 531 428 533 430
rect 527 427 533 428
rect 481 422 495 424
rect 480 420 495 422
rect 498 421 509 423
rect 480 418 481 420
rect 483 418 485 420
rect 480 416 485 418
rect 498 419 499 421
rect 501 419 509 421
rect 498 417 509 419
rect 481 411 485 416
rect 481 409 482 411
rect 484 409 485 411
rect 481 399 485 409
rect 488 406 489 412
rect 505 407 509 417
rect 529 407 533 427
rect 505 406 533 407
rect 505 405 518 406
rect 505 403 506 405
rect 508 404 518 405
rect 520 404 529 406
rect 531 404 533 406
rect 508 403 533 404
rect 505 401 509 403
rect 481 395 497 399
rect 493 394 506 395
rect 493 392 502 394
rect 504 392 506 394
rect 493 391 506 392
rect 295 384 301 385
rect 295 382 297 384
rect 299 382 301 384
rect 335 384 341 385
rect 335 382 337 384
rect 339 382 341 384
rect 370 384 374 386
rect 370 382 371 384
rect 373 382 374 384
rect 409 384 415 385
rect 409 382 411 384
rect 413 382 415 384
rect 444 384 448 386
rect 444 382 445 384
rect 447 382 448 384
rect 483 384 489 385
rect 483 382 485 384
rect 487 382 489 384
rect 518 384 522 386
rect 518 382 519 384
rect 521 382 522 384
rect -18 364 -16 366
rect -14 364 -12 366
rect -18 363 -12 364
rect -10 359 7 360
rect -10 357 3 359
rect 5 357 7 359
rect -10 356 7 357
rect 21 357 27 366
rect -25 345 -24 356
rect -10 352 -6 356
rect 21 355 23 357
rect 25 355 27 357
rect 21 354 27 355
rect 32 359 36 361
rect 32 357 33 359
rect 35 357 36 359
rect -21 348 -6 352
rect -21 335 -17 348
rect 32 352 36 357
rect 41 359 47 366
rect 70 364 71 366
rect 73 364 74 366
rect 41 357 43 359
rect 45 357 47 359
rect 41 356 47 357
rect 70 359 74 364
rect 70 357 71 359
rect 73 357 74 359
rect 70 355 74 357
rect 78 360 111 361
rect 78 358 107 360
rect 109 358 111 360
rect 78 357 111 358
rect 125 357 131 366
rect 32 351 33 352
rect 19 350 33 351
rect 35 350 36 352
rect 19 347 36 350
rect -2 339 4 340
rect -21 333 -20 335
rect -18 333 -17 335
rect -21 327 -17 333
rect -21 326 -3 327
rect -21 324 -7 326
rect -5 324 -3 326
rect -21 323 -3 324
rect 19 335 23 347
rect 78 346 82 357
rect 125 355 127 357
rect 129 355 131 357
rect 125 354 131 355
rect 136 359 140 361
rect 136 357 137 359
rect 139 357 140 359
rect 59 345 82 346
rect 59 343 61 345
rect 63 343 82 345
rect 59 342 82 343
rect 59 336 63 342
rect 19 333 20 335
rect 22 333 23 335
rect 19 328 23 333
rect 19 324 31 328
rect 15 321 16 323
rect 27 320 31 324
rect 52 332 63 336
rect 52 326 56 332
rect 78 336 82 342
rect 86 352 90 354
rect 86 350 87 352
rect 89 350 90 352
rect 86 345 90 350
rect 86 343 87 345
rect 89 344 90 345
rect 89 343 102 344
rect 86 340 102 343
rect 98 338 102 340
rect 98 336 103 338
rect 78 335 94 336
rect 78 333 90 335
rect 92 333 94 335
rect 78 332 94 333
rect 98 334 100 336
rect 102 334 103 336
rect 98 332 103 334
rect 52 324 53 326
rect 55 324 56 326
rect 52 322 56 324
rect 98 328 102 332
rect 78 324 102 328
rect 78 321 82 324
rect 27 319 47 320
rect 78 319 79 321
rect 81 319 82 321
rect 27 317 43 319
rect 45 317 47 319
rect 27 316 47 317
rect 65 318 71 319
rect 65 316 67 318
rect 69 316 71 318
rect 78 317 82 319
rect 136 352 140 357
rect 145 359 151 366
rect 174 364 175 366
rect 177 364 178 366
rect 145 357 147 359
rect 149 357 151 359
rect 145 356 151 357
rect 174 359 178 364
rect 174 357 175 359
rect 177 357 178 359
rect 174 355 178 357
rect 182 360 215 361
rect 182 358 211 360
rect 213 358 215 360
rect 182 357 215 358
rect 228 359 234 366
rect 228 357 230 359
rect 232 357 234 359
rect 136 351 137 352
rect 123 350 137 351
rect 139 350 140 352
rect 123 347 140 350
rect 123 335 127 347
rect 182 346 186 357
rect 228 356 234 357
rect 239 359 243 361
rect 239 357 240 359
rect 242 357 243 359
rect 163 345 186 346
rect 163 343 165 345
rect 167 343 186 345
rect 163 342 186 343
rect 163 336 167 342
rect 123 333 124 335
rect 126 333 127 335
rect 123 328 127 333
rect 123 324 135 328
rect 119 321 120 323
rect -18 313 -12 314
rect -18 311 -16 313
rect -14 311 -12 313
rect -18 310 -12 311
rect 1 313 7 314
rect 1 311 3 313
rect 5 311 7 313
rect 1 310 7 311
rect 65 310 71 316
rect 131 320 135 324
rect 156 332 167 336
rect 156 326 160 332
rect 182 336 186 342
rect 190 352 194 354
rect 190 350 191 352
rect 193 350 194 352
rect 190 345 194 350
rect 190 343 191 345
rect 193 344 194 345
rect 193 343 206 344
rect 190 340 206 343
rect 202 338 206 340
rect 202 336 207 338
rect 182 335 198 336
rect 182 333 194 335
rect 196 333 198 335
rect 182 332 198 333
rect 202 334 204 336
rect 206 334 207 336
rect 202 332 207 334
rect 156 324 157 326
rect 159 324 160 326
rect 156 322 160 324
rect 202 328 206 332
rect 182 324 206 328
rect 239 352 243 357
rect 248 357 254 366
rect 295 364 297 366
rect 299 364 301 366
rect 295 363 301 364
rect 335 364 337 366
rect 339 364 341 366
rect 335 363 341 364
rect 370 364 371 366
rect 373 364 374 366
rect 370 362 374 364
rect 409 364 411 366
rect 413 364 415 366
rect 409 363 415 364
rect 444 364 445 366
rect 447 364 448 366
rect 444 362 448 364
rect 483 364 485 366
rect 487 364 489 366
rect 483 363 489 364
rect 518 364 519 366
rect 521 364 522 366
rect 518 362 522 364
rect 248 355 250 357
rect 252 355 254 357
rect 276 359 293 360
rect 276 357 278 359
rect 280 357 293 359
rect 276 356 293 357
rect 248 354 254 355
rect 239 350 240 352
rect 242 351 243 352
rect 242 350 256 351
rect 239 347 256 350
rect 182 321 186 324
rect 131 319 151 320
rect 182 319 183 321
rect 185 319 186 321
rect 252 335 256 347
rect 252 333 253 335
rect 255 333 256 335
rect 252 328 256 333
rect 244 324 256 328
rect 289 352 293 356
rect 289 348 304 352
rect 279 339 285 340
rect 244 320 248 324
rect 259 321 260 323
rect 300 335 304 348
rect 307 345 308 356
rect 300 333 301 335
rect 303 333 304 335
rect 300 327 304 333
rect 286 326 304 327
rect 286 324 288 326
rect 290 324 304 326
rect 286 323 304 324
rect 345 356 358 357
rect 345 354 354 356
rect 356 354 358 356
rect 345 353 358 354
rect 333 349 349 353
rect 333 339 337 349
rect 419 356 432 357
rect 357 345 361 347
rect 333 337 334 339
rect 336 337 337 339
rect 333 332 337 337
rect 332 330 337 332
rect 357 343 358 345
rect 360 344 385 345
rect 360 343 370 344
rect 357 342 370 343
rect 372 342 381 344
rect 383 342 385 344
rect 357 341 385 342
rect 357 331 361 341
rect 332 328 333 330
rect 335 328 337 330
rect 350 329 361 331
rect 332 326 347 328
rect 333 324 347 326
rect 350 327 351 329
rect 353 327 361 329
rect 350 325 361 327
rect 131 317 147 319
rect 149 317 151 319
rect 131 316 151 317
rect 169 318 175 319
rect 169 316 171 318
rect 173 316 175 318
rect 182 317 186 319
rect 228 319 248 320
rect 228 317 230 319
rect 232 317 248 319
rect 228 316 248 317
rect 169 310 175 316
rect 336 318 340 320
rect 336 316 337 318
rect 339 316 340 318
rect 276 313 282 314
rect 276 311 278 313
rect 280 311 282 313
rect 276 310 282 311
rect 295 313 301 314
rect 295 311 297 313
rect 299 311 301 313
rect 295 310 301 311
rect 336 310 340 316
rect 343 319 347 324
rect 381 321 385 341
rect 369 320 375 321
rect 343 318 358 319
rect 343 316 354 318
rect 356 316 358 318
rect 343 315 358 316
rect 369 318 371 320
rect 373 318 375 320
rect 369 310 375 318
rect 379 320 385 321
rect 379 318 381 320
rect 383 318 385 320
rect 379 317 385 318
rect 419 354 428 356
rect 430 354 432 356
rect 419 353 432 354
rect 407 349 423 353
rect 407 339 411 349
rect 493 356 506 357
rect 431 345 435 347
rect 407 337 408 339
rect 410 337 411 339
rect 407 332 411 337
rect 431 343 432 345
rect 434 344 459 345
rect 434 343 444 344
rect 431 342 444 343
rect 446 342 455 344
rect 457 342 459 344
rect 431 341 459 342
rect 406 330 411 332
rect 431 331 435 341
rect 406 328 407 330
rect 409 328 411 330
rect 424 329 435 331
rect 406 326 421 328
rect 407 324 421 326
rect 424 327 425 329
rect 427 327 435 329
rect 424 325 435 327
rect 410 318 414 320
rect 410 316 411 318
rect 413 316 414 318
rect 410 310 414 316
rect 417 319 421 324
rect 455 321 459 341
rect 443 320 449 321
rect 417 318 432 319
rect 417 316 428 318
rect 430 316 432 318
rect 417 315 432 316
rect 443 318 445 320
rect 447 318 449 320
rect 443 310 449 318
rect 453 320 459 321
rect 453 318 455 320
rect 457 318 459 320
rect 453 317 459 318
rect 493 354 502 356
rect 504 354 506 356
rect 493 353 506 354
rect 481 349 497 353
rect 481 339 485 349
rect 505 345 509 347
rect 481 337 482 339
rect 484 337 485 339
rect 481 332 485 337
rect 488 336 489 342
rect 505 343 506 345
rect 508 344 533 345
rect 508 343 518 344
rect 505 342 518 343
rect 520 342 529 344
rect 531 342 533 344
rect 505 341 533 342
rect 480 330 485 332
rect 505 331 509 341
rect 480 328 481 330
rect 483 328 485 330
rect 498 329 509 331
rect 480 326 495 328
rect 481 324 495 326
rect 498 327 499 329
rect 501 327 509 329
rect 498 325 509 327
rect 484 318 488 320
rect 484 316 485 318
rect 487 316 488 318
rect 484 310 488 316
rect 491 319 495 324
rect 529 321 533 341
rect 517 320 523 321
rect 491 318 506 319
rect 491 316 502 318
rect 504 316 506 318
rect 491 315 506 316
rect 517 318 519 320
rect 521 318 523 320
rect 517 310 523 318
rect 527 320 533 321
rect 527 318 529 320
rect 531 318 533 320
rect 527 317 533 318
rect -18 293 -12 294
rect -18 291 -16 293
rect -14 291 -12 293
rect -18 290 -12 291
rect 1 293 7 294
rect 1 291 3 293
rect 5 291 7 293
rect 1 290 7 291
rect 65 288 71 294
rect 27 287 47 288
rect 27 285 43 287
rect 45 285 47 287
rect 65 286 67 288
rect 69 286 71 288
rect 65 285 71 286
rect 78 285 82 287
rect 27 284 47 285
rect -21 280 -3 281
rect -21 278 -7 280
rect -5 278 -3 280
rect -21 277 -3 278
rect -21 271 -17 277
rect -21 269 -20 271
rect -18 269 -17 271
rect -25 248 -24 259
rect -21 256 -17 269
rect -2 264 4 265
rect -21 252 -6 256
rect -10 248 -6 252
rect 15 281 16 283
rect 27 280 31 284
rect 78 283 79 285
rect 81 283 82 285
rect 19 276 31 280
rect 19 271 23 276
rect 19 269 20 271
rect 22 269 23 271
rect 19 257 23 269
rect 52 280 56 282
rect 52 278 53 280
rect 55 278 56 280
rect 52 272 56 278
rect 78 280 82 283
rect 78 276 102 280
rect 52 268 63 272
rect 19 254 36 257
rect 19 253 33 254
rect 32 252 33 253
rect 35 252 36 254
rect 21 249 27 250
rect -10 247 7 248
rect -10 245 3 247
rect 5 245 7 247
rect -10 244 7 245
rect 21 247 23 249
rect 25 247 27 249
rect -18 240 -12 241
rect -18 238 -16 240
rect -14 238 -12 240
rect 21 238 27 247
rect 32 247 36 252
rect 59 262 63 268
rect 98 272 102 276
rect 78 271 94 272
rect 78 269 90 271
rect 92 269 94 271
rect 78 268 94 269
rect 98 270 103 272
rect 98 268 100 270
rect 102 268 103 270
rect 78 262 82 268
rect 98 266 103 268
rect 98 264 102 266
rect 59 261 82 262
rect 59 259 61 261
rect 63 259 82 261
rect 59 258 82 259
rect 32 245 33 247
rect 35 245 36 247
rect 32 243 36 245
rect 41 247 47 248
rect 41 245 43 247
rect 45 245 47 247
rect 41 238 47 245
rect 70 247 74 249
rect 70 245 71 247
rect 73 245 74 247
rect 70 240 74 245
rect 78 247 82 258
rect 86 261 102 264
rect 86 259 87 261
rect 89 260 102 261
rect 89 259 90 260
rect 86 254 90 259
rect 86 252 87 254
rect 89 252 90 254
rect 86 250 90 252
rect 169 288 175 294
rect 276 293 282 294
rect 276 291 278 293
rect 280 291 282 293
rect 276 290 282 291
rect 295 293 301 294
rect 295 291 297 293
rect 299 291 301 293
rect 295 290 301 291
rect 131 287 151 288
rect 131 285 147 287
rect 149 285 151 287
rect 169 286 171 288
rect 173 286 175 288
rect 169 285 175 286
rect 182 285 186 287
rect 131 284 151 285
rect 119 281 120 283
rect 131 280 135 284
rect 182 283 183 285
rect 185 283 186 285
rect 228 287 248 288
rect 228 285 230 287
rect 232 285 248 287
rect 228 284 248 285
rect 123 276 135 280
rect 123 271 127 276
rect 123 269 124 271
rect 126 269 127 271
rect 123 257 127 269
rect 156 280 160 282
rect 156 278 157 280
rect 159 278 160 280
rect 156 272 160 278
rect 182 280 186 283
rect 182 276 206 280
rect 156 268 167 272
rect 123 254 140 257
rect 123 253 137 254
rect 136 252 137 253
rect 139 252 140 254
rect 125 249 131 250
rect 125 247 127 249
rect 129 247 131 249
rect 78 246 111 247
rect 78 244 107 246
rect 109 244 111 246
rect 78 243 111 244
rect 70 238 71 240
rect 73 238 74 240
rect 125 238 131 247
rect 136 247 140 252
rect 163 262 167 268
rect 202 272 206 276
rect 182 271 198 272
rect 182 269 194 271
rect 196 269 198 271
rect 182 268 198 269
rect 202 270 207 272
rect 202 268 204 270
rect 206 268 207 270
rect 182 262 186 268
rect 202 266 207 268
rect 202 264 206 266
rect 163 261 186 262
rect 163 259 165 261
rect 167 259 186 261
rect 163 258 186 259
rect 136 245 137 247
rect 139 245 140 247
rect 136 243 140 245
rect 145 247 151 248
rect 145 245 147 247
rect 149 245 151 247
rect 145 238 151 245
rect 174 247 178 249
rect 174 245 175 247
rect 177 245 178 247
rect 174 240 178 245
rect 182 247 186 258
rect 190 261 206 264
rect 190 259 191 261
rect 193 260 206 261
rect 193 259 194 260
rect 190 254 194 259
rect 244 280 248 284
rect 259 281 260 283
rect 244 276 256 280
rect 252 271 256 276
rect 252 269 253 271
rect 255 269 256 271
rect 190 252 191 254
rect 193 252 194 254
rect 190 250 194 252
rect 252 257 256 269
rect 336 288 340 294
rect 336 286 337 288
rect 339 286 340 288
rect 336 284 340 286
rect 343 288 358 289
rect 343 286 354 288
rect 356 286 358 288
rect 343 285 358 286
rect 369 286 375 294
rect 410 288 414 294
rect 286 280 304 281
rect 286 278 288 280
rect 290 278 304 280
rect 286 277 304 278
rect 300 271 304 277
rect 300 269 301 271
rect 303 269 304 271
rect 279 264 285 265
rect 239 254 256 257
rect 239 252 240 254
rect 242 253 256 254
rect 242 252 243 253
rect 228 247 234 248
rect 182 246 215 247
rect 182 244 211 246
rect 213 244 215 246
rect 182 243 215 244
rect 228 245 230 247
rect 232 245 234 247
rect 174 238 175 240
rect 177 238 178 240
rect 228 238 234 245
rect 239 247 243 252
rect 300 256 304 269
rect 289 252 304 256
rect 239 245 240 247
rect 242 245 243 247
rect 239 243 243 245
rect 248 249 254 250
rect 248 247 250 249
rect 252 247 254 249
rect 289 248 293 252
rect 307 248 308 259
rect 248 238 254 247
rect 276 247 293 248
rect 276 245 278 247
rect 280 245 293 247
rect 276 244 293 245
rect 343 280 347 285
rect 369 284 371 286
rect 373 284 375 286
rect 369 283 375 284
rect 379 286 385 287
rect 379 284 381 286
rect 383 284 385 286
rect 379 283 385 284
rect 333 278 347 280
rect 332 276 347 278
rect 350 277 361 279
rect 332 274 333 276
rect 335 274 337 276
rect 332 272 337 274
rect 350 275 351 277
rect 353 275 361 277
rect 350 273 361 275
rect 333 267 337 272
rect 333 265 334 267
rect 336 265 337 267
rect 333 255 337 265
rect 357 263 361 273
rect 381 263 385 283
rect 357 262 385 263
rect 357 261 370 262
rect 357 259 358 261
rect 360 260 370 261
rect 372 260 381 262
rect 383 260 385 262
rect 360 259 385 260
rect 410 286 411 288
rect 413 286 414 288
rect 410 284 414 286
rect 417 288 432 289
rect 417 286 428 288
rect 430 286 432 288
rect 417 285 432 286
rect 443 286 449 294
rect 484 288 488 294
rect 417 280 421 285
rect 443 284 445 286
rect 447 284 449 286
rect 443 283 449 284
rect 453 286 459 287
rect 453 284 455 286
rect 457 284 459 286
rect 453 283 459 284
rect 407 278 421 280
rect 406 276 421 278
rect 424 277 435 279
rect 406 274 407 276
rect 409 274 411 276
rect 406 272 411 274
rect 424 275 425 277
rect 427 275 435 277
rect 424 273 435 275
rect 357 257 361 259
rect 333 251 349 255
rect 345 250 358 251
rect 345 248 354 250
rect 356 248 358 250
rect 345 247 358 248
rect 407 267 411 272
rect 407 265 408 267
rect 410 265 411 267
rect 407 255 411 265
rect 431 263 435 273
rect 455 263 459 283
rect 431 262 459 263
rect 431 261 444 262
rect 431 259 432 261
rect 434 260 444 261
rect 446 260 455 262
rect 457 260 459 262
rect 434 259 459 260
rect 484 286 485 288
rect 487 286 488 288
rect 484 284 488 286
rect 491 288 506 289
rect 491 286 502 288
rect 504 286 506 288
rect 491 285 506 286
rect 517 286 523 294
rect 431 257 435 259
rect 407 251 423 255
rect 419 250 432 251
rect 419 248 428 250
rect 430 248 432 250
rect 419 247 432 248
rect 491 280 495 285
rect 517 284 519 286
rect 521 284 523 286
rect 517 283 523 284
rect 527 286 533 287
rect 527 284 529 286
rect 531 284 533 286
rect 527 283 533 284
rect 481 278 495 280
rect 480 276 495 278
rect 498 277 509 279
rect 480 274 481 276
rect 483 274 485 276
rect 480 272 485 274
rect 498 275 499 277
rect 501 275 509 277
rect 498 273 509 275
rect 481 267 485 272
rect 481 265 482 267
rect 484 265 485 267
rect 481 255 485 265
rect 488 262 489 268
rect 505 263 509 273
rect 529 263 533 283
rect 505 262 533 263
rect 505 261 518 262
rect 505 259 506 261
rect 508 260 518 261
rect 520 260 529 262
rect 531 260 533 262
rect 508 259 533 260
rect 505 257 509 259
rect 481 251 497 255
rect 493 250 506 251
rect 493 248 502 250
rect 504 248 506 250
rect 493 247 506 248
rect 295 240 301 241
rect 295 238 297 240
rect 299 238 301 240
rect 335 240 341 241
rect 335 238 337 240
rect 339 238 341 240
rect 370 240 374 242
rect 370 238 371 240
rect 373 238 374 240
rect 409 240 415 241
rect 409 238 411 240
rect 413 238 415 240
rect 444 240 448 242
rect 444 238 445 240
rect 447 238 448 240
rect 483 240 489 241
rect 483 238 485 240
rect 487 238 489 240
rect 518 240 522 242
rect 518 238 519 240
rect 521 238 522 240
rect -18 220 -16 222
rect -14 220 -12 222
rect -18 219 -12 220
rect -10 215 7 216
rect -10 213 3 215
rect 5 213 7 215
rect -10 212 7 213
rect 21 213 27 222
rect -25 201 -24 212
rect -10 208 -6 212
rect 21 211 23 213
rect 25 211 27 213
rect 21 210 27 211
rect 32 215 36 217
rect 32 213 33 215
rect 35 213 36 215
rect -21 204 -6 208
rect -21 191 -17 204
rect 32 208 36 213
rect 41 215 47 222
rect 70 220 71 222
rect 73 220 74 222
rect 41 213 43 215
rect 45 213 47 215
rect 41 212 47 213
rect 70 215 74 220
rect 70 213 71 215
rect 73 213 74 215
rect 70 211 74 213
rect 78 216 111 217
rect 78 214 107 216
rect 109 214 111 216
rect 78 213 111 214
rect 125 213 131 222
rect 32 207 33 208
rect 19 206 33 207
rect 35 206 36 208
rect 19 203 36 206
rect -2 195 4 196
rect -21 189 -20 191
rect -18 189 -17 191
rect -21 183 -17 189
rect -21 182 -3 183
rect -21 180 -7 182
rect -5 180 -3 182
rect -21 179 -3 180
rect 19 191 23 203
rect 78 202 82 213
rect 125 211 127 213
rect 129 211 131 213
rect 125 210 131 211
rect 136 215 140 217
rect 136 213 137 215
rect 139 213 140 215
rect 59 201 82 202
rect 59 199 61 201
rect 63 199 82 201
rect 59 198 82 199
rect 59 192 63 198
rect 19 189 20 191
rect 22 189 23 191
rect 19 184 23 189
rect 19 180 31 184
rect 15 177 16 179
rect 27 176 31 180
rect 52 188 63 192
rect 52 182 56 188
rect 78 192 82 198
rect 86 208 90 210
rect 86 206 87 208
rect 89 206 90 208
rect 86 201 90 206
rect 86 199 87 201
rect 89 200 90 201
rect 89 199 102 200
rect 86 196 102 199
rect 98 194 102 196
rect 98 192 103 194
rect 78 191 94 192
rect 78 189 90 191
rect 92 189 94 191
rect 78 188 94 189
rect 98 190 100 192
rect 102 190 103 192
rect 98 188 103 190
rect 52 180 53 182
rect 55 180 56 182
rect 52 178 56 180
rect 98 184 102 188
rect 78 180 102 184
rect 78 177 82 180
rect 27 175 47 176
rect 78 175 79 177
rect 81 175 82 177
rect 27 173 43 175
rect 45 173 47 175
rect 27 172 47 173
rect 65 174 71 175
rect 65 172 67 174
rect 69 172 71 174
rect 78 173 82 175
rect 136 208 140 213
rect 145 215 151 222
rect 174 220 175 222
rect 177 220 178 222
rect 145 213 147 215
rect 149 213 151 215
rect 145 212 151 213
rect 174 215 178 220
rect 174 213 175 215
rect 177 213 178 215
rect 174 211 178 213
rect 182 216 215 217
rect 182 214 211 216
rect 213 214 215 216
rect 182 213 215 214
rect 228 215 234 222
rect 228 213 230 215
rect 232 213 234 215
rect 136 207 137 208
rect 123 206 137 207
rect 139 206 140 208
rect 123 203 140 206
rect 123 191 127 203
rect 182 202 186 213
rect 228 212 234 213
rect 239 215 243 217
rect 239 213 240 215
rect 242 213 243 215
rect 163 201 186 202
rect 163 199 165 201
rect 167 199 186 201
rect 163 198 186 199
rect 163 192 167 198
rect 123 189 124 191
rect 126 189 127 191
rect 123 184 127 189
rect 123 180 135 184
rect 119 177 120 179
rect -18 169 -12 170
rect -18 167 -16 169
rect -14 167 -12 169
rect -18 166 -12 167
rect 1 169 7 170
rect 1 167 3 169
rect 5 167 7 169
rect 1 166 7 167
rect 65 166 71 172
rect 131 176 135 180
rect 156 188 167 192
rect 156 182 160 188
rect 182 192 186 198
rect 190 208 194 210
rect 190 206 191 208
rect 193 206 194 208
rect 190 201 194 206
rect 190 199 191 201
rect 193 200 194 201
rect 193 199 206 200
rect 190 196 206 199
rect 202 194 206 196
rect 202 192 207 194
rect 182 191 198 192
rect 182 189 194 191
rect 196 189 198 191
rect 182 188 198 189
rect 202 190 204 192
rect 206 190 207 192
rect 202 188 207 190
rect 156 180 157 182
rect 159 180 160 182
rect 156 178 160 180
rect 202 184 206 188
rect 182 180 206 184
rect 239 208 243 213
rect 248 213 254 222
rect 295 220 297 222
rect 299 220 301 222
rect 295 219 301 220
rect 335 220 337 222
rect 339 220 341 222
rect 335 219 341 220
rect 370 220 371 222
rect 373 220 374 222
rect 370 218 374 220
rect 409 220 411 222
rect 413 220 415 222
rect 409 219 415 220
rect 444 220 445 222
rect 447 220 448 222
rect 444 218 448 220
rect 483 220 485 222
rect 487 220 489 222
rect 483 219 489 220
rect 518 220 519 222
rect 521 220 522 222
rect 518 218 522 220
rect 248 211 250 213
rect 252 211 254 213
rect 276 215 293 216
rect 276 213 278 215
rect 280 213 293 215
rect 276 212 293 213
rect 248 210 254 211
rect 239 206 240 208
rect 242 207 243 208
rect 242 206 256 207
rect 239 203 256 206
rect 182 177 186 180
rect 131 175 151 176
rect 182 175 183 177
rect 185 175 186 177
rect 252 191 256 203
rect 252 189 253 191
rect 255 189 256 191
rect 252 184 256 189
rect 244 180 256 184
rect 289 208 293 212
rect 289 204 304 208
rect 279 195 285 196
rect 244 176 248 180
rect 259 177 260 179
rect 300 191 304 204
rect 307 201 308 212
rect 300 189 301 191
rect 303 189 304 191
rect 300 183 304 189
rect 286 182 304 183
rect 286 180 288 182
rect 290 180 304 182
rect 286 179 304 180
rect 345 212 358 213
rect 345 210 354 212
rect 356 210 358 212
rect 345 209 358 210
rect 333 205 349 209
rect 333 195 337 205
rect 419 212 432 213
rect 357 201 361 203
rect 333 193 334 195
rect 336 193 337 195
rect 333 188 337 193
rect 332 186 337 188
rect 357 199 358 201
rect 360 200 385 201
rect 360 199 370 200
rect 357 198 370 199
rect 372 198 381 200
rect 383 198 385 200
rect 357 197 385 198
rect 357 187 361 197
rect 332 184 333 186
rect 335 184 337 186
rect 350 185 361 187
rect 332 182 347 184
rect 333 180 347 182
rect 350 183 351 185
rect 353 183 361 185
rect 350 181 361 183
rect 131 173 147 175
rect 149 173 151 175
rect 131 172 151 173
rect 169 174 175 175
rect 169 172 171 174
rect 173 172 175 174
rect 182 173 186 175
rect 228 175 248 176
rect 228 173 230 175
rect 232 173 248 175
rect 228 172 248 173
rect 169 166 175 172
rect 336 174 340 176
rect 336 172 337 174
rect 339 172 340 174
rect 276 169 282 170
rect 276 167 278 169
rect 280 167 282 169
rect 276 166 282 167
rect 295 169 301 170
rect 295 167 297 169
rect 299 167 301 169
rect 295 166 301 167
rect 336 166 340 172
rect 343 175 347 180
rect 381 177 385 197
rect 369 176 375 177
rect 343 174 358 175
rect 343 172 354 174
rect 356 172 358 174
rect 343 171 358 172
rect 369 174 371 176
rect 373 174 375 176
rect 369 166 375 174
rect 379 176 385 177
rect 379 174 381 176
rect 383 174 385 176
rect 379 173 385 174
rect 419 210 428 212
rect 430 210 432 212
rect 419 209 432 210
rect 407 205 423 209
rect 407 195 411 205
rect 493 212 506 213
rect 431 201 435 203
rect 407 193 408 195
rect 410 193 411 195
rect 407 188 411 193
rect 431 199 432 201
rect 434 200 459 201
rect 434 199 444 200
rect 431 198 444 199
rect 446 198 455 200
rect 457 198 459 200
rect 431 197 459 198
rect 406 186 411 188
rect 431 187 435 197
rect 406 184 407 186
rect 409 184 411 186
rect 424 185 435 187
rect 406 182 421 184
rect 407 180 421 182
rect 424 183 425 185
rect 427 183 435 185
rect 424 181 435 183
rect 410 174 414 176
rect 410 172 411 174
rect 413 172 414 174
rect 410 166 414 172
rect 417 175 421 180
rect 455 177 459 197
rect 443 176 449 177
rect 417 174 432 175
rect 417 172 428 174
rect 430 172 432 174
rect 417 171 432 172
rect 443 174 445 176
rect 447 174 449 176
rect 443 166 449 174
rect 453 176 459 177
rect 453 174 455 176
rect 457 174 459 176
rect 453 173 459 174
rect 493 210 502 212
rect 504 210 506 212
rect 493 209 506 210
rect 481 205 497 209
rect 481 195 485 205
rect 505 201 509 203
rect 481 193 482 195
rect 484 193 485 195
rect 481 188 485 193
rect 488 192 489 198
rect 505 199 506 201
rect 508 200 533 201
rect 508 199 518 200
rect 505 198 518 199
rect 520 198 529 200
rect 531 198 533 200
rect 505 197 533 198
rect 480 186 485 188
rect 505 187 509 197
rect 480 184 481 186
rect 483 184 485 186
rect 498 185 509 187
rect 480 182 495 184
rect 481 180 495 182
rect 498 183 499 185
rect 501 183 509 185
rect 498 181 509 183
rect 484 174 488 176
rect 484 172 485 174
rect 487 172 488 174
rect 484 166 488 172
rect 491 175 495 180
rect 529 177 533 197
rect 517 176 523 177
rect 491 174 506 175
rect 491 172 502 174
rect 504 172 506 174
rect 491 171 506 172
rect 517 174 519 176
rect 521 174 523 176
rect 517 166 523 174
rect 527 176 533 177
rect 527 174 529 176
rect 531 174 533 176
rect 527 173 533 174
<< via1 >>
rect 4 413 6 415
rect 4 400 6 402
rect 36 422 38 424
rect 12 400 14 402
rect 61 422 63 424
rect 69 422 71 424
rect 44 398 46 400
rect 53 398 55 400
rect 108 405 110 407
rect 116 413 118 415
rect 140 422 142 424
rect 131 413 133 415
rect 165 422 167 424
rect 139 405 141 407
rect 148 398 150 400
rect 212 417 214 419
rect 157 398 159 400
rect 237 422 239 424
rect 229 405 231 407
rect 277 422 279 424
rect 261 408 263 410
rect 277 405 279 407
rect 309 407 311 409
rect 326 415 328 417
rect 341 405 343 407
rect 368 415 370 417
rect 400 411 402 413
rect 417 413 419 415
rect 490 411 492 413
rect 516 420 518 422
rect -28 358 -26 360
rect 4 346 6 348
rect 12 346 14 348
rect 44 348 46 350
rect 4 333 6 335
rect 53 348 55 350
rect 36 324 38 326
rect 108 341 110 343
rect 61 324 63 326
rect 148 348 150 350
rect 116 333 118 335
rect 139 341 141 343
rect 157 348 159 350
rect 131 333 133 335
rect 140 324 142 326
rect 165 324 167 326
rect 229 341 231 343
rect 212 329 214 331
rect 236 324 238 326
rect 277 341 279 343
rect 261 338 263 340
rect 309 339 311 341
rect 277 324 279 326
rect 326 331 328 333
rect 341 341 343 343
rect 368 331 370 333
rect 400 335 402 337
rect 417 333 419 335
rect 490 335 492 337
rect 516 326 518 328
rect -36 273 -34 275
rect 4 269 6 271
rect 4 256 6 258
rect 36 278 38 280
rect 12 256 14 258
rect 61 278 63 280
rect 69 278 71 280
rect 44 254 46 256
rect 53 254 55 256
rect 108 261 110 263
rect 116 269 118 271
rect 140 278 142 280
rect 131 269 133 271
rect 165 278 167 280
rect 139 261 141 263
rect 148 254 150 256
rect 212 273 214 275
rect 157 254 159 256
rect 237 278 239 280
rect 229 261 231 263
rect 277 278 279 280
rect 261 264 263 266
rect 277 261 279 263
rect 309 263 311 265
rect 326 271 328 273
rect 341 261 343 263
rect 368 271 370 273
rect 400 267 402 269
rect 417 269 419 271
rect 490 267 492 269
rect 516 276 518 278
rect -28 214 -26 216
rect 4 202 6 204
rect 12 202 14 204
rect 44 204 46 206
rect 4 189 6 191
rect 53 204 55 206
rect 36 180 38 182
rect 108 197 110 199
rect 61 180 63 182
rect 148 204 150 206
rect 116 189 118 191
rect 139 197 141 199
rect 157 204 159 206
rect 140 180 142 182
rect 165 180 167 182
rect 229 197 231 199
rect 212 185 214 187
rect 236 180 238 182
rect 277 197 279 199
rect 261 194 263 196
rect 309 195 311 197
rect 277 180 279 182
rect 326 187 328 189
rect 341 197 343 199
rect 368 187 370 189
rect 400 191 402 193
rect 417 189 419 191
rect 490 191 492 193
rect 516 182 518 184
<< via2 >>
rect 69 422 71 424
rect 237 422 239 424
rect 277 422 279 424
rect 131 413 133 415
rect 53 398 55 400
rect 229 405 231 407
rect 277 405 279 407
rect -28 358 -26 360
rect 53 348 55 350
rect 131 333 133 335
rect 229 341 231 343
rect 277 341 279 343
rect 61 324 63 326
rect 236 324 238 326
rect 277 324 279 326
rect 69 278 71 280
rect 237 278 239 280
rect 277 278 279 280
rect -36 273 -34 275
rect 131 269 133 271
rect 53 254 55 256
rect 229 261 231 263
rect 277 261 279 263
rect -28 214 -26 216
rect 53 204 55 206
rect 229 197 231 199
rect 277 197 279 199
rect 61 180 63 182
rect 236 180 238 182
rect 277 180 279 182
<< labels >>
rlabel polyct1 382 210 382 210 1 s0
rlabel polyct1 456 210 456 210 1 s0
rlabel polyct1 530 210 530 210 1 s1
rlabel alu1 383 227 383 227 1 vdd!
rlabel alu1 501 161 501 161 1 vss!
rlabel polyct1 382 250 382 250 5 s0
rlabel polyct1 456 250 456 250 5 s0
rlabel polyct1 530 250 530 250 5 s1
rlabel alu1 383 233 383 233 5 vdd!
rlabel alu1 501 299 501 299 5 vss!
rlabel polyct1 382 354 382 354 1 s0
rlabel polyct1 456 354 456 354 1 s0
rlabel polyct1 530 354 530 354 1 s1
rlabel alu1 383 371 383 371 1 vdd!
rlabel alu1 501 305 501 305 1 vss!
rlabel polyct1 382 394 382 394 5 s0
rlabel polyct1 456 394 456 394 5 s0
rlabel polyct1 530 394 530 394 5 s1
rlabel alu1 383 377 383 377 5 vdd!
rlabel alu1 501 443 501 443 5 vss!
rlabel pwell 211 328 215 332 1 sum2
rlabel alu1 473 336 477 340 1 aluout2
rlabel alu1 473 407 477 410 1 aluout3
rlabel pwell 211 416 215 420 1 sum3
rlabel alu1 -27 418 -27 418 1 cout
rlabel alu1 37 418 37 418 1 a3
rlabel alu2 48 325 48 325 1 a2
rlabel alu2 49 399 49 399 1 b3
rlabel alu2 49 349 49 349 1 b2
rlabel alu2 49 255 49 255 1 b1
rlabel alu1 37 274 37 274 1 a1
rlabel pwell 211 272 215 276 1 sum1
rlabel alu1 473 263 477 266 1 aluout1
rlabel alu2 48 181 48 181 1 a0
rlabel alu2 49 205 49 205 1 b0
rlabel pwell 211 184 215 188 1 sum0
rlabel alu1 473 192 477 196 1 aluout0
rlabel alu1 141 187 141 187 1 cin
<< end >>
