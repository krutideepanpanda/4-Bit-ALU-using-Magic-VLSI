* SPICE3 file created from ALU1bit.ext - technology: scmos

.option scale=0.055u

M1000 zn a vdd vdd pmos w=13 l=2
+  ad=104 pd=42 as=2950 ps=900
M1001 an_1 cin vdd vdd pmos w=18 l=2
+  ad=144 pd=52 as=0 ps=0
M1002 vdd a_266_32# a_220_80# vdd pmos w=19 l=2
+  ad=0 pd=0 as=342 ps=112
M1003 vdd zn co vdd pmos w=18 l=2
+  ad=0 pd=0 as=116 ps=50
M1004 vdd b bn vdd pmos w=27 l=2
+  ad=0 pd=0 as=294 ps=136
M1005 a_n103_34# cin vss vss nmos w=11 l=2
+  ad=55 pd=32 as=2057 ps=802
M1006 i1 a_8_19# vss vss nmos w=19 l=2
+  ad=152 pd=54 as=0 ps=0
M1007 vss cmd0 a_266_32# vss nmos w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1008 vss co zn_2 vss nmos w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1009 an_1 cin vss vss nmos w=9 l=2
+  ad=72 pd=34 as=0 ps=0
M1010 vss cmd0 a_220_16# vss nmos w=12 l=2
+  ad=0 pd=0 as=246 ps=94
M1011 s bn an vdd pmos w=18 l=2
+  ad=189 pd=70 as=144 ps=52
M1012 vdd zn_2 a_n269_41# vdd pmos w=18 l=2
+  ad=0 pd=0 as=126 ps=50
M1013 zn_1 cin vdd vdd pmos w=13 l=2
+  ad=104 pd=42 as=0 ps=0
M1014 a_230_16# i2 a_220_16# vss nmos w=12 l=2
+  ad=120 pd=44 as=0 ps=0
M1015 a_8_19# a vdd vdd pmos w=20 l=2
+  ad=203 pd=62 as=0 ps=0
M1016 s b an vss nmos w=9 l=2
+  ad=87 pd=40 as=72 ps=34
M1017 vdd zn_1 c1 vdd pmos w=18 l=2
+  ad=0 pd=0 as=116 ps=50
M1018 vdd s zn_1 vdd pmos w=13 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 vss b bn vss nmos w=9 l=2
+  ad=0 pd=0 as=57 ps=32
M1020 i2 a_108_60# vdd vdd pmos w=39 l=2
+  ad=312 pd=94 as=0 ps=0
M1021 a_220_80# i1 a_254_80# vdd pmos w=19 l=2
+  ad=0 pd=0 as=114 ps=50
M1022 vss b a_18_19# vss nmos w=18 l=2
+  ad=0 pd=0 as=244 ps=76
M1023 zn_1 s a_n103_34# vss nmos w=11 l=2
+  ad=67 pd=36 as=0 ps=0
M1024 vss an_1 a_n40_30# vss nmos w=12 l=2
+  ad=0 pd=0 as=60 ps=34
M1025 zn_2 c1 vss vss nmos w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1026 vss zn co vss nmos w=9 l=2
+  ad=0 pd=0 as=57 ps=32
M1027 an a vdd vdd pmos w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 i1 a_8_19# vdd vdd pmos w=39 l=2
+  ad=312 pd=94 as=0 ps=0
M1029 vss b a_108_60# vss nmos w=10 l=2
+  ad=0 pd=0 as=103 ps=42
M1030 bn_1 an_1 i0 vdd pmos w=27 l=2
+  ad=294 pd=136 as=189 ps=70
M1031 a_n40_30# bn_1 i0 vss nmos w=12 l=2
+  ad=0 pd=0 as=87 ps=40
M1032 a_254_80# a_218_34# nq vdd pmos w=19 l=2
+  ad=0 pd=0 as=388 ps=128
M1033 an a vss vss nmos w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 a_220_16# i1 a_254_16# vss nmos w=12 l=2
+  ad=0 pd=0 as=72 ps=36
M1035 vdd b a_122_61# vdd pmos w=29 l=2
+  ad=0 pd=0 as=174 ps=70
M1036 vss zn_2 a_n269_41# vss nmos w=9 l=2
+  ad=0 pd=0 as=57 ps=32
M1037 vss zn_1 c1 vss nmos w=9 l=2
+  ad=0 pd=0 as=57 ps=32
M1038 nq i0 a_286_80# vdd pmos w=19 l=2
+  ad=0 pd=0 as=114 ps=50
M1039 vdd b zn vdd pmos w=13 l=2
+  ad=0 pd=0 as=0 ps=0
M1040 vdd s bn_1 vdd pmos w=27 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 a_254_16# cmd1 nq vss nmos w=12 l=2
+  ad=0 pd=0 as=300 ps=112
M1042 a_218_34# cmd1 vdd vdd pmos w=14 l=2
+  ad=112 pd=44 as=0 ps=0
M1043 a_108_60# a vss vss nmos w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1044 nq i0 a_286_12# vss nmos w=12 l=2
+  ad=0 pd=0 as=72 ps=36
M1045 i0 bn_1 an_1 vdd pmos w=18 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 a_122_61# a a_108_60# vdd pmos w=29 l=2
+  ad=0 pd=0 as=354 ps=84
M1047 nq cmd1 a_230_80# vdd pmos w=18 l=2
+  ad=0 pd=0 as=185 ps=58
M1048 zn b a_n207_34# vss nmos w=11 l=2
+  ad=67 pd=36 as=55 ps=32
M1049 vss an a_n144_30# vss nmos w=12 l=2
+  ad=0 pd=0 as=60 ps=34
M1050 a_286_80# cmd0 vdd vdd pmos w=19 l=2
+  ad=0 pd=0 as=0 ps=0
M1051 zn_2 co a_n247_66# vdd pmos w=21 l=2
+  ad=117 pd=56 as=105 ps=52
M1052 a_18_19# a a_8_19# vss nmos w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1053 vdd cmd0 a_266_32# vdd pmos w=14 l=2
+  ad=0 pd=0 as=112 ps=44
M1054 i0 s an_1 vss nmos w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 bn an s vdd pmos w=27 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 a_n207_34# a vss vss nmos w=11 l=2
+  ad=0 pd=0 as=0 ps=0
M1057 a_n144_30# bn s vss nmos w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1058 a_n247_66# c1 vdd vdd pmos w=21 l=2
+  ad=0 pd=0 as=0 ps=0
M1059 a_286_12# a_266_32# vss vss nmos w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 vss s bn_1 vss nmos w=9 l=2
+  ad=0 pd=0 as=57 ps=32
M1061 i2 a_108_60# vss vss nmos w=19 l=2
+  ad=152 pd=54 as=0 ps=0
M1062 nq a_218_34# a_230_16# vss nmos w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1063 vdd b a_8_19# vdd pmos w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 a_230_80# i2 a_220_80# vdd pmos w=19 l=2
+  ad=0 pd=0 as=0 ps=0
M1065 a_218_34# cmd1 vss vss nmos w=8 l=2
+  ad=64 pd=32 as=0 ps=0
