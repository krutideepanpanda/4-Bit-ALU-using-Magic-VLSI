magic
tech scmos
timestamp 1636283722
<< ab >>
rect 44 302 50 307
rect 148 302 154 307
rect -31 301 217 302
rect -31 300 131 301
rect -31 297 -14 300
rect -10 297 27 300
rect -31 296 27 297
rect 31 299 131 300
rect 31 296 80 299
rect 82 297 131 299
rect 135 299 217 301
rect 135 297 183 299
rect 82 296 183 297
rect 187 296 217 299
rect -31 270 217 296
rect -31 238 49 270
rect 50 238 153 270
rect 154 238 217 270
rect -31 236 217 238
rect -31 232 -14 236
rect -9 232 26 236
rect 30 232 79 236
rect 83 232 130 236
rect 134 232 183 236
rect 187 232 217 236
rect -31 228 217 232
rect -31 224 -14 228
rect -9 224 26 228
rect 30 224 79 228
rect 83 224 130 228
rect 134 224 183 228
rect 187 224 217 228
rect -31 222 217 224
rect -31 190 49 222
rect 50 190 153 222
rect 154 190 217 222
rect -31 164 217 190
rect -31 163 27 164
rect -31 160 -14 163
rect -10 160 27 163
rect 31 161 80 164
rect 82 163 183 164
rect 82 161 131 163
rect 31 160 131 161
rect -31 159 131 160
rect 135 161 183 163
rect 187 161 217 164
rect 135 159 217 161
rect -31 157 217 159
rect -31 156 131 157
rect -31 153 -14 156
rect -10 153 27 156
rect -31 152 27 153
rect 31 155 131 156
rect 31 152 80 155
rect 82 153 131 155
rect 135 155 217 157
rect 135 153 183 155
rect 82 152 183 153
rect 187 152 217 155
rect -31 148 217 152
rect -37 144 217 148
rect -31 134 217 144
rect -37 130 217 134
rect -31 126 217 130
rect -31 94 49 126
rect 50 94 153 126
rect 154 94 217 126
rect -31 92 217 94
rect -31 88 -14 92
rect -9 88 26 92
rect 30 88 79 92
rect 83 88 130 92
rect 134 88 183 92
rect 187 88 217 92
rect -31 84 217 88
rect -31 80 -14 84
rect -9 80 26 84
rect 30 80 79 84
rect 83 80 130 84
rect 134 80 183 84
rect 187 80 217 84
rect -31 78 217 80
rect -31 77 49 78
rect -31 72 -29 77
rect -25 72 49 77
rect -31 57 49 72
rect -32 53 49 57
rect -29 49 49 53
rect -31 46 49 49
rect 50 46 153 78
rect 154 46 217 78
rect -31 20 217 46
rect -31 19 27 20
rect -31 16 -14 19
rect -10 16 27 19
rect 31 17 80 20
rect 82 19 183 20
rect 82 17 131 19
rect 31 16 131 17
rect -31 15 131 16
rect 135 17 183 19
rect 187 17 217 20
rect 135 15 217 17
rect -31 14 217 15
rect 226 300 266 302
rect 226 296 244 300
rect 248 296 266 300
rect 226 287 266 296
rect 226 285 237 287
rect 239 285 253 287
rect 255 285 266 287
rect 226 271 266 285
rect 226 269 261 271
rect 263 269 266 271
rect 226 268 266 269
rect 226 266 253 268
rect 255 266 266 268
rect 226 251 266 266
rect 226 249 240 251
rect 242 249 266 251
rect 226 236 266 249
rect 226 232 244 236
rect 248 232 266 236
rect 226 228 266 232
rect 226 224 244 228
rect 248 224 266 228
rect 226 211 266 224
rect 226 209 240 211
rect 242 209 266 211
rect 226 194 266 209
rect 226 192 253 194
rect 255 192 266 194
rect 226 191 266 192
rect 226 189 261 191
rect 263 189 266 191
rect 226 175 266 189
rect 226 173 237 175
rect 239 173 253 175
rect 255 173 266 175
rect 226 164 266 173
rect 226 160 244 164
rect 248 160 266 164
rect 226 156 266 160
rect 226 152 244 156
rect 248 152 266 156
rect 226 143 266 152
rect 226 141 237 143
rect 239 141 253 143
rect 255 141 266 143
rect 226 127 266 141
rect 226 125 261 127
rect 263 125 266 127
rect 226 124 266 125
rect 226 122 253 124
rect 255 122 266 124
rect 226 107 266 122
rect 226 105 240 107
rect 242 105 266 107
rect 226 92 266 105
rect 226 88 244 92
rect 248 88 266 92
rect 226 84 266 88
rect 226 80 244 84
rect 248 80 266 84
rect 226 67 266 80
rect 226 65 240 67
rect 242 65 266 67
rect 226 50 266 65
rect 226 48 253 50
rect 255 48 266 50
rect 226 47 266 48
rect 226 45 261 47
rect 263 45 266 47
rect 226 31 266 45
rect 226 29 237 31
rect 239 29 253 31
rect 255 29 266 31
rect 226 20 266 29
rect 226 16 244 20
rect 248 16 266 20
rect 226 14 266 16
rect 274 300 314 302
rect 274 297 292 300
rect 296 297 314 300
rect 274 280 314 297
rect 274 278 294 280
rect 296 278 314 280
rect 274 268 314 278
rect 274 266 301 268
rect 303 266 314 268
rect 274 263 314 266
rect 274 261 309 263
rect 311 261 314 263
rect 274 247 314 261
rect 274 245 284 247
rect 286 245 301 247
rect 303 245 314 247
rect 274 236 314 245
rect 274 232 292 236
rect 296 232 314 236
rect 274 228 314 232
rect 274 224 292 228
rect 296 224 314 228
rect 274 215 314 224
rect 274 213 284 215
rect 286 213 301 215
rect 303 213 314 215
rect 274 199 314 213
rect 274 197 309 199
rect 311 197 314 199
rect 274 194 314 197
rect 274 192 301 194
rect 303 192 314 194
rect 274 182 314 192
rect 274 180 294 182
rect 296 180 314 182
rect 274 163 314 180
rect 274 160 292 163
rect 296 160 314 163
rect 274 156 314 160
rect 274 153 292 156
rect 296 153 314 156
rect 274 136 314 153
rect 274 134 294 136
rect 296 134 314 136
rect 274 124 314 134
rect 274 122 301 124
rect 303 122 314 124
rect 274 119 314 122
rect 274 117 309 119
rect 311 117 314 119
rect 274 103 314 117
rect 274 101 284 103
rect 286 101 301 103
rect 303 101 314 103
rect 274 92 314 101
rect 274 88 292 92
rect 296 88 314 92
rect 274 84 314 88
rect 274 80 292 84
rect 296 80 314 84
rect 274 71 314 80
rect 274 69 284 71
rect 286 69 301 71
rect 303 69 314 71
rect 274 55 314 69
rect 274 53 309 55
rect 311 53 314 55
rect 274 50 314 53
rect 274 48 301 50
rect 303 48 314 50
rect 274 38 314 48
rect 274 36 294 38
rect 296 36 314 38
rect 274 19 314 36
rect 274 16 292 19
rect 296 16 314 19
rect 274 14 314 16
rect 323 299 387 302
rect 323 297 354 299
rect 356 297 387 299
rect 323 289 387 297
rect 323 285 349 289
rect 351 285 387 289
rect 323 279 387 285
rect 323 277 374 279
rect 376 277 387 279
rect 323 275 354 277
rect 356 275 387 277
rect 323 274 387 275
rect 323 272 382 274
rect 384 272 387 274
rect 323 271 387 272
rect 323 269 326 271
rect 328 269 366 271
rect 370 269 387 271
rect 323 267 358 269
rect 360 267 387 269
rect 323 265 334 267
rect 336 265 342 267
rect 344 265 387 267
rect 323 263 387 265
rect 323 261 350 263
rect 352 262 387 263
rect 352 261 370 262
rect 323 260 370 261
rect 372 260 387 262
rect 323 255 387 260
rect 323 253 374 255
rect 376 253 387 255
rect 323 251 387 253
rect 323 248 349 251
rect 353 248 387 251
rect 323 247 387 248
rect 323 245 334 247
rect 336 245 382 247
rect 384 245 387 247
rect 323 235 387 245
rect 323 233 354 235
rect 356 233 387 235
rect 323 227 387 233
rect 323 225 354 227
rect 356 225 387 227
rect 323 215 387 225
rect 323 213 334 215
rect 336 213 382 215
rect 384 213 387 215
rect 323 212 387 213
rect 323 209 349 212
rect 353 209 387 212
rect 323 207 387 209
rect 323 205 374 207
rect 376 205 387 207
rect 323 200 387 205
rect 323 199 370 200
rect 323 197 350 199
rect 352 198 370 199
rect 372 198 387 200
rect 352 197 387 198
rect 323 195 387 197
rect 323 193 334 195
rect 336 193 342 195
rect 344 193 387 195
rect 323 191 358 193
rect 360 191 387 193
rect 323 189 326 191
rect 328 189 366 191
rect 370 189 387 191
rect 323 188 387 189
rect 323 186 382 188
rect 384 186 387 188
rect 323 185 387 186
rect 323 183 354 185
rect 356 183 387 185
rect 323 181 374 183
rect 376 181 387 183
rect 323 175 387 181
rect 323 171 349 175
rect 351 171 387 175
rect 323 163 387 171
rect 323 161 354 163
rect 356 161 387 163
rect 323 155 387 161
rect 323 153 354 155
rect 356 153 387 155
rect 323 145 387 153
rect 323 141 349 145
rect 351 141 387 145
rect 323 135 387 141
rect 323 133 374 135
rect 376 133 387 135
rect 323 131 354 133
rect 356 131 387 133
rect 323 130 387 131
rect 323 128 382 130
rect 384 128 387 130
rect 323 127 387 128
rect 323 125 326 127
rect 328 125 366 127
rect 370 125 387 127
rect 323 123 358 125
rect 360 123 387 125
rect 323 121 334 123
rect 336 121 342 123
rect 344 121 387 123
rect 323 119 387 121
rect 323 117 350 119
rect 352 118 387 119
rect 352 117 370 118
rect 323 116 370 117
rect 372 116 387 118
rect 323 111 387 116
rect 323 109 374 111
rect 376 109 387 111
rect 323 107 387 109
rect 323 104 349 107
rect 353 104 387 107
rect 323 103 387 104
rect 323 101 334 103
rect 336 101 382 103
rect 384 101 387 103
rect 323 91 387 101
rect 323 89 354 91
rect 356 89 387 91
rect 323 83 387 89
rect 323 81 354 83
rect 356 81 387 83
rect 323 71 387 81
rect 323 69 334 71
rect 336 69 382 71
rect 384 69 387 71
rect 323 68 387 69
rect 323 65 349 68
rect 353 65 387 68
rect 323 63 387 65
rect 323 61 374 63
rect 376 61 387 63
rect 323 56 387 61
rect 323 55 370 56
rect 323 53 350 55
rect 352 54 370 55
rect 372 54 387 56
rect 352 53 387 54
rect 323 51 387 53
rect 323 49 334 51
rect 336 49 342 51
rect 344 49 387 51
rect 323 47 358 49
rect 360 47 387 49
rect 323 45 326 47
rect 328 45 366 47
rect 370 45 387 47
rect 323 44 387 45
rect 323 42 382 44
rect 384 42 387 44
rect 323 41 387 42
rect 323 39 354 41
rect 356 39 387 41
rect 323 37 374 39
rect 376 37 387 39
rect 323 31 387 37
rect 323 27 349 31
rect 351 27 387 31
rect 323 19 387 27
rect 323 17 354 19
rect 356 17 387 19
rect 323 14 387 17
rect 397 299 461 302
rect 397 297 428 299
rect 430 297 461 299
rect 397 289 461 297
rect 397 285 423 289
rect 425 285 461 289
rect 397 279 461 285
rect 397 277 448 279
rect 450 277 461 279
rect 397 275 428 277
rect 430 275 461 277
rect 397 274 461 275
rect 397 272 456 274
rect 458 272 461 274
rect 397 271 461 272
rect 397 269 400 271
rect 402 269 440 271
rect 442 269 461 271
rect 397 267 432 269
rect 434 267 461 269
rect 397 265 408 267
rect 410 265 416 267
rect 418 265 461 267
rect 397 263 461 265
rect 397 261 424 263
rect 426 262 461 263
rect 426 261 444 262
rect 397 260 444 261
rect 446 260 461 262
rect 397 255 461 260
rect 397 253 448 255
rect 450 253 461 255
rect 397 251 461 253
rect 397 248 423 251
rect 427 248 461 251
rect 397 247 461 248
rect 397 245 408 247
rect 410 245 456 247
rect 458 245 461 247
rect 397 235 461 245
rect 397 233 428 235
rect 430 233 461 235
rect 397 227 461 233
rect 397 225 428 227
rect 430 225 461 227
rect 397 215 461 225
rect 397 213 408 215
rect 410 213 456 215
rect 458 213 461 215
rect 397 212 461 213
rect 397 209 423 212
rect 427 209 461 212
rect 397 207 461 209
rect 397 205 448 207
rect 450 205 461 207
rect 397 200 461 205
rect 397 199 444 200
rect 397 197 424 199
rect 426 198 444 199
rect 446 198 461 200
rect 426 197 461 198
rect 397 195 461 197
rect 397 193 408 195
rect 410 193 416 195
rect 418 193 461 195
rect 397 191 432 193
rect 434 191 461 193
rect 397 189 400 191
rect 402 189 440 191
rect 442 189 461 191
rect 397 188 461 189
rect 397 186 456 188
rect 458 186 461 188
rect 397 185 461 186
rect 397 183 428 185
rect 430 183 461 185
rect 397 181 448 183
rect 450 181 461 183
rect 397 175 461 181
rect 397 171 423 175
rect 425 171 461 175
rect 397 163 461 171
rect 397 161 428 163
rect 430 161 461 163
rect 397 155 461 161
rect 397 153 428 155
rect 430 153 461 155
rect 397 145 461 153
rect 397 141 423 145
rect 425 141 461 145
rect 397 135 461 141
rect 397 133 448 135
rect 450 133 461 135
rect 397 131 428 133
rect 430 131 461 133
rect 397 130 461 131
rect 397 128 456 130
rect 458 128 461 130
rect 397 127 461 128
rect 397 125 400 127
rect 402 125 440 127
rect 442 125 461 127
rect 397 123 432 125
rect 434 123 461 125
rect 397 121 408 123
rect 410 121 416 123
rect 418 121 461 123
rect 397 119 461 121
rect 397 117 424 119
rect 426 118 461 119
rect 426 117 444 118
rect 397 116 444 117
rect 446 116 461 118
rect 397 111 461 116
rect 397 109 448 111
rect 450 109 461 111
rect 397 107 461 109
rect 397 104 423 107
rect 427 104 461 107
rect 397 103 461 104
rect 397 101 408 103
rect 410 101 456 103
rect 458 101 461 103
rect 397 91 461 101
rect 397 89 428 91
rect 430 89 461 91
rect 397 83 461 89
rect 397 81 428 83
rect 430 81 461 83
rect 397 71 461 81
rect 397 69 408 71
rect 410 69 456 71
rect 458 69 461 71
rect 397 68 461 69
rect 397 65 423 68
rect 427 65 461 68
rect 397 63 461 65
rect 397 61 448 63
rect 450 61 461 63
rect 397 56 461 61
rect 397 55 444 56
rect 397 53 424 55
rect 426 54 444 55
rect 446 54 461 56
rect 426 53 461 54
rect 397 51 461 53
rect 397 49 408 51
rect 410 49 416 51
rect 418 49 461 51
rect 397 47 432 49
rect 434 47 461 49
rect 397 45 400 47
rect 402 45 440 47
rect 442 45 461 47
rect 397 44 461 45
rect 397 42 456 44
rect 458 42 461 44
rect 397 41 461 42
rect 397 39 428 41
rect 430 39 461 41
rect 397 37 448 39
rect 450 37 461 39
rect 397 31 461 37
rect 397 27 423 31
rect 425 27 461 31
rect 397 19 461 27
rect 397 17 428 19
rect 430 17 461 19
rect 397 14 461 17
rect 471 299 535 302
rect 471 297 502 299
rect 504 297 535 299
rect 471 289 535 297
rect 471 285 497 289
rect 499 285 535 289
rect 471 279 535 285
rect 471 277 522 279
rect 524 277 535 279
rect 471 275 502 277
rect 504 275 535 277
rect 471 274 535 275
rect 471 272 530 274
rect 532 272 535 274
rect 471 271 535 272
rect 471 269 474 271
rect 476 269 514 271
rect 516 269 535 271
rect 471 268 506 269
rect 471 266 474 268
rect 476 267 506 268
rect 508 267 535 269
rect 476 266 482 267
rect 471 265 482 266
rect 484 265 490 267
rect 492 265 535 267
rect 471 263 535 265
rect 471 261 498 263
rect 500 262 535 263
rect 500 261 518 262
rect 471 260 518 261
rect 520 260 535 262
rect 471 255 535 260
rect 471 253 522 255
rect 524 253 535 255
rect 471 251 535 253
rect 471 248 497 251
rect 501 248 535 251
rect 471 247 535 248
rect 471 245 482 247
rect 484 245 530 247
rect 532 245 535 247
rect 471 235 535 245
rect 471 233 502 235
rect 504 233 535 235
rect 471 227 535 233
rect 471 225 502 227
rect 504 225 535 227
rect 471 215 535 225
rect 471 213 482 215
rect 484 213 530 215
rect 532 213 535 215
rect 471 212 535 213
rect 471 209 497 212
rect 501 209 535 212
rect 471 207 535 209
rect 471 205 522 207
rect 524 205 535 207
rect 471 200 535 205
rect 471 199 518 200
rect 471 197 498 199
rect 500 198 518 199
rect 520 198 535 200
rect 500 197 535 198
rect 471 195 535 197
rect 471 194 482 195
rect 471 192 474 194
rect 476 193 482 194
rect 484 193 490 195
rect 492 193 535 195
rect 476 192 506 193
rect 471 191 506 192
rect 508 191 535 193
rect 471 189 474 191
rect 476 189 514 191
rect 516 189 535 191
rect 471 188 535 189
rect 471 186 530 188
rect 532 186 535 188
rect 471 185 535 186
rect 471 183 502 185
rect 504 183 535 185
rect 471 181 522 183
rect 524 181 535 183
rect 471 175 535 181
rect 471 171 497 175
rect 499 171 535 175
rect 471 163 535 171
rect 471 161 502 163
rect 504 161 535 163
rect 471 155 535 161
rect 471 153 502 155
rect 504 153 535 155
rect 471 145 535 153
rect 471 141 497 145
rect 499 141 535 145
rect 471 135 535 141
rect 471 133 522 135
rect 524 133 535 135
rect 471 131 502 133
rect 504 131 535 133
rect 471 130 535 131
rect 471 128 530 130
rect 532 128 535 130
rect 471 127 535 128
rect 471 125 474 127
rect 476 125 514 127
rect 516 125 535 127
rect 471 124 506 125
rect 471 122 474 124
rect 476 123 506 124
rect 508 123 535 125
rect 476 122 482 123
rect 471 121 482 122
rect 484 121 490 123
rect 492 121 535 123
rect 471 119 535 121
rect 471 117 498 119
rect 500 118 535 119
rect 500 117 518 118
rect 471 116 518 117
rect 520 116 535 118
rect 471 111 535 116
rect 471 109 522 111
rect 524 109 535 111
rect 471 107 535 109
rect 471 104 497 107
rect 501 104 535 107
rect 471 103 535 104
rect 471 101 482 103
rect 484 101 530 103
rect 532 101 535 103
rect 471 91 535 101
rect 471 89 502 91
rect 504 89 535 91
rect 471 83 535 89
rect 471 81 502 83
rect 504 81 535 83
rect 471 71 535 81
rect 471 69 482 71
rect 484 69 530 71
rect 532 69 535 71
rect 471 68 535 69
rect 471 65 497 68
rect 501 65 535 68
rect 471 63 535 65
rect 471 61 522 63
rect 524 61 535 63
rect 471 56 535 61
rect 471 55 518 56
rect 471 53 498 55
rect 500 54 518 55
rect 520 54 535 56
rect 500 53 535 54
rect 471 51 535 53
rect 471 50 482 51
rect 471 48 474 50
rect 476 49 482 50
rect 484 49 490 51
rect 492 49 535 51
rect 476 48 506 49
rect 471 47 506 48
rect 508 47 535 49
rect 471 45 474 47
rect 476 45 514 47
rect 516 45 535 47
rect 471 44 535 45
rect 471 42 530 44
rect 532 42 535 44
rect 471 41 535 42
rect 471 39 502 41
rect 504 39 535 41
rect 471 37 522 39
rect 524 37 535 39
rect 471 31 535 37
rect 471 27 497 31
rect 499 27 535 31
rect 471 19 535 27
rect 471 17 502 19
rect 504 17 535 19
rect 471 14 535 17
rect 44 9 50 14
rect 148 9 154 14
<< nwell >>
rect -37 190 540 270
rect -37 46 540 126
<< pwell >>
rect -37 270 540 307
rect -37 126 540 190
rect -37 9 540 46
<< poly >>
rect -22 285 -20 290
rect -12 282 -10 287
rect -2 282 0 287
rect 18 287 20 291
rect 31 289 33 294
rect 38 289 40 294
rect 61 298 86 300
rect 61 290 63 298
rect 74 290 76 294
rect 84 290 86 298
rect 94 293 96 298
rect 101 293 103 298
rect 58 288 63 290
rect 58 285 60 288
rect -22 273 -20 276
rect -12 273 -10 276
rect -22 271 -16 273
rect -22 269 -20 271
rect -18 269 -16 271
rect -22 267 -16 269
rect -12 271 -6 273
rect -12 269 -10 271
rect -8 269 -6 271
rect -12 267 -6 269
rect -22 264 -20 267
rect -9 257 -7 267
rect -2 266 0 276
rect 18 273 20 278
rect 31 273 33 278
rect 18 271 24 273
rect 18 269 20 271
rect 22 269 24 271
rect 18 267 24 269
rect 28 271 34 273
rect 28 269 30 271
rect 32 269 34 271
rect 28 267 34 269
rect -2 264 4 266
rect -2 262 0 264
rect 2 262 4 264
rect 18 263 20 267
rect -2 260 4 262
rect -2 257 0 260
rect -22 241 -20 246
rect 28 256 30 267
rect 38 265 40 278
rect 122 287 124 291
rect 135 289 137 294
rect 142 289 144 294
rect 165 298 190 300
rect 165 290 167 298
rect 178 290 180 294
rect 188 290 190 298
rect 198 293 200 298
rect 205 293 207 298
rect 74 278 76 281
rect 67 276 76 278
rect 84 277 86 281
rect 94 278 96 281
rect 58 268 60 276
rect 67 274 69 276
rect 71 274 76 276
rect 67 272 76 274
rect 92 276 96 278
rect 92 273 94 276
rect 74 268 76 272
rect 88 271 94 273
rect 101 272 103 281
rect 162 288 167 290
rect 162 285 164 288
rect 122 273 124 278
rect 135 273 137 278
rect 88 269 90 271
rect 92 269 94 271
rect 55 266 68 268
rect 74 266 84 268
rect 88 267 94 269
rect 55 265 57 266
rect 38 263 44 265
rect 38 261 40 263
rect 42 261 44 263
rect 38 259 44 261
rect 51 263 57 265
rect 66 263 68 266
rect 82 263 84 266
rect 92 263 94 267
rect 98 270 104 272
rect 98 268 100 270
rect 102 268 104 270
rect 98 266 104 268
rect 102 263 104 266
rect 122 271 128 273
rect 122 269 124 271
rect 126 269 128 271
rect 122 267 128 269
rect 132 271 138 273
rect 132 269 134 271
rect 136 269 138 271
rect 132 267 138 269
rect 122 263 124 267
rect 51 261 53 263
rect 55 261 57 263
rect 51 259 57 261
rect 38 256 40 259
rect 18 241 20 245
rect 28 238 30 243
rect 38 238 40 243
rect -9 232 -7 236
rect -2 232 0 236
rect 82 241 84 245
rect 92 241 94 245
rect 66 232 68 236
rect 132 256 134 267
rect 142 265 144 278
rect 235 289 237 294
rect 242 289 244 294
rect 359 298 378 300
rect 178 278 180 281
rect 171 276 180 278
rect 188 277 190 281
rect 198 278 200 281
rect 162 268 164 276
rect 171 274 173 276
rect 175 274 180 276
rect 171 272 180 274
rect 196 276 200 278
rect 196 273 198 276
rect 178 268 180 272
rect 192 271 198 273
rect 205 272 207 281
rect 255 287 257 291
rect 332 290 334 295
rect 342 290 344 295
rect 349 290 351 295
rect 359 290 361 298
rect 366 290 368 294
rect 283 282 285 287
rect 293 282 295 287
rect 303 285 305 290
rect 192 269 194 271
rect 196 269 198 271
rect 159 266 172 268
rect 178 266 188 268
rect 192 267 198 269
rect 159 265 161 266
rect 142 263 148 265
rect 142 261 144 263
rect 146 261 148 263
rect 142 259 148 261
rect 155 263 161 265
rect 170 263 172 266
rect 186 263 188 266
rect 196 263 198 267
rect 202 270 208 272
rect 202 268 204 270
rect 206 268 208 270
rect 202 266 208 268
rect 206 263 208 266
rect 235 265 237 278
rect 242 273 244 278
rect 255 273 257 278
rect 376 288 378 298
rect 433 298 452 300
rect 406 290 408 295
rect 416 290 418 295
rect 423 290 425 295
rect 433 290 435 298
rect 440 290 442 294
rect 332 278 334 281
rect 331 276 337 278
rect 241 271 247 273
rect 241 269 243 271
rect 245 269 247 271
rect 241 267 247 269
rect 251 271 257 273
rect 251 269 253 271
rect 255 269 257 271
rect 251 267 257 269
rect 231 263 237 265
rect 155 261 157 263
rect 159 261 161 263
rect 155 259 161 261
rect 142 256 144 259
rect 122 241 124 245
rect 132 238 134 243
rect 142 238 144 243
rect 102 232 104 236
rect 186 241 188 245
rect 196 241 198 245
rect 170 232 172 236
rect 231 261 233 263
rect 235 261 237 263
rect 231 259 237 261
rect 235 256 237 259
rect 245 256 247 267
rect 255 263 257 267
rect 283 266 285 276
rect 293 273 295 276
rect 303 273 305 276
rect 289 271 295 273
rect 289 269 291 271
rect 293 269 295 271
rect 289 267 295 269
rect 299 271 305 273
rect 331 274 333 276
rect 335 274 337 276
rect 331 272 337 274
rect 299 269 301 271
rect 303 269 305 271
rect 299 267 305 269
rect 279 264 285 266
rect 279 262 281 264
rect 283 262 285 264
rect 279 260 285 262
rect 283 257 285 260
rect 290 257 292 267
rect 303 264 305 267
rect 235 238 237 243
rect 245 238 247 243
rect 255 241 257 245
rect 206 232 208 236
rect 332 254 334 272
rect 342 268 344 282
rect 349 279 351 282
rect 349 277 355 279
rect 349 275 351 277
rect 353 275 355 277
rect 349 273 355 275
rect 359 269 361 282
rect 339 266 345 268
rect 339 264 341 266
rect 343 264 345 266
rect 339 262 345 264
rect 349 267 361 269
rect 366 278 368 282
rect 366 276 372 278
rect 366 274 368 276
rect 370 274 372 276
rect 366 267 372 274
rect 303 241 305 246
rect 283 232 285 236
rect 290 232 292 236
rect 342 252 344 262
rect 349 252 351 267
rect 356 261 362 263
rect 356 259 358 261
rect 360 259 362 261
rect 356 257 362 259
rect 359 252 361 257
rect 366 252 368 267
rect 376 264 378 282
rect 450 288 452 298
rect 507 298 526 300
rect 480 290 482 295
rect 490 290 492 295
rect 497 290 499 295
rect 507 290 509 298
rect 514 290 516 294
rect 406 278 408 281
rect 405 276 411 278
rect 405 274 407 276
rect 409 274 411 276
rect 405 272 411 274
rect 376 253 378 256
rect 406 254 408 272
rect 416 268 418 282
rect 423 279 425 282
rect 423 277 429 279
rect 423 275 425 277
rect 427 275 429 277
rect 423 273 429 275
rect 433 269 435 282
rect 413 266 419 268
rect 413 264 415 266
rect 417 264 419 266
rect 413 262 419 264
rect 423 267 435 269
rect 440 273 442 282
rect 440 271 446 273
rect 440 269 442 271
rect 444 269 446 271
rect 440 267 446 269
rect 376 251 385 253
rect 379 249 381 251
rect 383 249 385 251
rect 379 247 385 249
rect 416 252 418 262
rect 423 252 425 267
rect 430 261 436 263
rect 430 259 432 261
rect 434 259 436 261
rect 430 257 436 259
rect 433 252 435 257
rect 440 252 442 267
rect 450 264 452 282
rect 524 288 526 298
rect 480 278 482 281
rect 479 276 485 278
rect 479 274 481 276
rect 483 274 485 276
rect 479 272 485 274
rect 450 253 452 256
rect 480 254 482 272
rect 490 268 492 282
rect 497 279 499 282
rect 497 277 503 279
rect 497 275 499 277
rect 501 275 503 277
rect 497 273 503 275
rect 507 269 509 282
rect 487 266 493 268
rect 487 264 489 266
rect 491 264 493 266
rect 487 262 493 264
rect 497 267 509 269
rect 514 273 516 282
rect 514 271 520 273
rect 514 269 516 271
rect 518 269 520 271
rect 514 267 520 269
rect 450 251 459 253
rect 453 249 455 251
rect 457 249 459 251
rect 453 247 459 249
rect 490 252 492 262
rect 497 252 499 267
rect 504 261 510 263
rect 504 259 506 261
rect 508 259 510 261
rect 504 257 510 259
rect 507 252 509 257
rect 514 252 516 267
rect 524 264 526 282
rect 524 253 526 256
rect 524 251 533 253
rect 527 249 529 251
rect 531 249 533 251
rect 527 247 533 249
rect 332 232 334 236
rect 342 232 344 236
rect 349 232 351 236
rect 359 232 361 236
rect 366 232 368 236
rect 406 232 408 236
rect 416 232 418 236
rect 423 232 425 236
rect 433 232 435 236
rect 440 232 442 236
rect 480 232 482 236
rect 490 232 492 236
rect 497 232 499 236
rect 507 232 509 236
rect 514 232 516 236
rect -9 224 -7 228
rect -2 224 0 228
rect -22 214 -20 219
rect 66 224 68 228
rect 18 215 20 219
rect 28 217 30 222
rect 38 217 40 222
rect -22 193 -20 196
rect -9 193 -7 203
rect -2 200 0 203
rect -2 198 4 200
rect -2 196 0 198
rect 2 196 4 198
rect -2 194 4 196
rect -22 191 -16 193
rect -22 189 -20 191
rect -18 189 -16 191
rect -22 187 -16 189
rect -12 191 -6 193
rect -12 189 -10 191
rect -8 189 -6 191
rect -12 187 -6 189
rect -22 184 -20 187
rect -12 184 -10 187
rect -2 184 0 194
rect 18 193 20 197
rect 28 193 30 204
rect 38 201 40 204
rect 38 199 44 201
rect 38 197 40 199
rect 42 197 44 199
rect 38 195 44 197
rect 51 199 57 201
rect 51 197 53 199
rect 55 197 57 199
rect 102 224 104 228
rect 82 215 84 219
rect 92 215 94 219
rect 170 224 172 228
rect 122 215 124 219
rect 132 217 134 222
rect 142 217 144 222
rect 51 195 57 197
rect 18 191 24 193
rect 18 189 20 191
rect 22 189 24 191
rect 18 187 24 189
rect 28 191 34 193
rect 28 189 30 191
rect 32 189 34 191
rect 28 187 34 189
rect 18 182 20 187
rect 31 182 33 187
rect 38 182 40 195
rect 55 194 57 195
rect 66 194 68 197
rect 82 194 84 197
rect 55 192 68 194
rect 74 192 84 194
rect 92 193 94 197
rect 102 194 104 197
rect 58 184 60 192
rect 74 188 76 192
rect 67 186 76 188
rect 88 191 94 193
rect 88 189 90 191
rect 92 189 94 191
rect 88 187 94 189
rect 98 192 104 194
rect 98 190 100 192
rect 102 190 104 192
rect 98 188 104 190
rect 122 193 124 197
rect 132 193 134 204
rect 142 201 144 204
rect 142 199 148 201
rect 142 197 144 199
rect 146 197 148 199
rect 142 195 148 197
rect 155 199 161 201
rect 155 197 157 199
rect 159 197 161 199
rect 206 224 208 228
rect 186 215 188 219
rect 196 215 198 219
rect 283 224 285 228
rect 290 224 292 228
rect 235 217 237 222
rect 245 217 247 222
rect 255 215 257 219
rect 235 201 237 204
rect 231 199 237 201
rect 231 197 233 199
rect 235 197 237 199
rect 155 195 161 197
rect 122 191 128 193
rect 122 189 124 191
rect 126 189 128 191
rect 67 184 69 186
rect 71 184 76 186
rect -22 170 -20 175
rect -12 173 -10 178
rect -2 173 0 178
rect 18 169 20 173
rect 67 182 76 184
rect 92 184 94 187
rect 74 179 76 182
rect 84 179 86 183
rect 92 182 96 184
rect 94 179 96 182
rect 101 179 103 188
rect 122 187 128 189
rect 132 191 138 193
rect 132 189 134 191
rect 136 189 138 191
rect 132 187 138 189
rect 122 182 124 187
rect 135 182 137 187
rect 142 182 144 195
rect 159 194 161 195
rect 170 194 172 197
rect 186 194 188 197
rect 159 192 172 194
rect 178 192 188 194
rect 196 193 198 197
rect 206 194 208 197
rect 231 195 237 197
rect 162 184 164 192
rect 178 188 180 192
rect 171 186 180 188
rect 192 191 198 193
rect 192 189 194 191
rect 196 189 198 191
rect 192 187 198 189
rect 202 192 208 194
rect 202 190 204 192
rect 206 190 208 192
rect 202 188 208 190
rect 171 184 173 186
rect 175 184 180 186
rect 58 172 60 175
rect 31 166 33 171
rect 38 166 40 171
rect 58 170 63 172
rect 61 162 63 170
rect 74 166 76 170
rect 84 162 86 170
rect 122 169 124 173
rect 171 182 180 184
rect 196 184 198 187
rect 178 179 180 182
rect 188 179 190 183
rect 196 182 200 184
rect 198 179 200 182
rect 205 179 207 188
rect 235 182 237 195
rect 245 193 247 204
rect 332 224 334 228
rect 342 224 344 228
rect 349 224 351 228
rect 359 224 361 228
rect 366 224 368 228
rect 406 224 408 228
rect 416 224 418 228
rect 423 224 425 228
rect 433 224 435 228
rect 440 224 442 228
rect 480 224 482 228
rect 490 224 492 228
rect 497 224 499 228
rect 507 224 509 228
rect 514 224 516 228
rect 303 214 305 219
rect 283 200 285 203
rect 279 198 285 200
rect 255 193 257 197
rect 279 196 281 198
rect 283 196 285 198
rect 279 194 285 196
rect 241 191 247 193
rect 241 189 243 191
rect 245 189 247 191
rect 241 187 247 189
rect 251 191 257 193
rect 251 189 253 191
rect 255 189 257 191
rect 251 187 257 189
rect 242 182 244 187
rect 255 182 257 187
rect 283 184 285 194
rect 290 193 292 203
rect 379 211 385 213
rect 379 209 381 211
rect 383 209 385 211
rect 303 193 305 196
rect 289 191 295 193
rect 289 189 291 191
rect 293 189 295 191
rect 289 187 295 189
rect 299 191 305 193
rect 299 189 301 191
rect 303 189 305 191
rect 299 187 305 189
rect 332 188 334 206
rect 342 198 344 208
rect 339 196 345 198
rect 339 194 341 196
rect 343 194 345 196
rect 339 192 345 194
rect 349 193 351 208
rect 359 203 361 208
rect 356 201 362 203
rect 356 199 358 201
rect 360 199 362 201
rect 356 197 362 199
rect 366 193 368 208
rect 376 207 385 209
rect 376 204 378 207
rect 453 211 459 213
rect 453 209 455 211
rect 457 209 459 211
rect 293 184 295 187
rect 303 184 305 187
rect 331 186 337 188
rect 331 184 333 186
rect 335 184 337 186
rect 162 172 164 175
rect 94 162 96 167
rect 101 162 103 167
rect 61 160 86 162
rect 135 166 137 171
rect 142 166 144 171
rect 162 170 167 172
rect 165 162 167 170
rect 178 166 180 170
rect 188 162 190 170
rect 198 162 200 167
rect 205 162 207 167
rect 235 166 237 171
rect 242 166 244 171
rect 165 160 190 162
rect 255 169 257 173
rect 283 173 285 178
rect 293 173 295 178
rect 331 182 337 184
rect 332 179 334 182
rect 303 170 305 175
rect 342 178 344 192
rect 349 191 361 193
rect 349 185 355 187
rect 349 183 351 185
rect 353 183 355 185
rect 349 181 355 183
rect 349 178 351 181
rect 359 178 361 191
rect 366 186 372 193
rect 366 184 368 186
rect 370 184 372 186
rect 366 182 372 184
rect 366 178 368 182
rect 376 178 378 196
rect 406 188 408 206
rect 416 198 418 208
rect 413 196 419 198
rect 413 194 415 196
rect 417 194 419 196
rect 413 192 419 194
rect 423 193 425 208
rect 433 203 435 208
rect 430 201 436 203
rect 430 199 432 201
rect 434 199 436 201
rect 430 197 436 199
rect 440 193 442 208
rect 450 207 459 209
rect 450 204 452 207
rect 527 211 533 213
rect 527 209 529 211
rect 531 209 533 211
rect 405 186 411 188
rect 405 184 407 186
rect 409 184 411 186
rect 405 182 411 184
rect 406 179 408 182
rect 332 165 334 170
rect 342 165 344 170
rect 349 165 351 170
rect 359 162 361 170
rect 366 166 368 170
rect 376 162 378 172
rect 416 178 418 192
rect 423 191 435 193
rect 423 185 429 187
rect 423 183 425 185
rect 427 183 429 185
rect 423 181 429 183
rect 423 178 425 181
rect 433 178 435 191
rect 440 191 446 193
rect 440 189 442 191
rect 444 189 446 191
rect 440 187 446 189
rect 440 178 442 187
rect 450 178 452 196
rect 480 188 482 206
rect 490 198 492 208
rect 487 196 493 198
rect 487 194 489 196
rect 491 194 493 196
rect 487 192 493 194
rect 497 193 499 208
rect 507 203 509 208
rect 504 201 510 203
rect 504 199 506 201
rect 508 199 510 201
rect 504 197 510 199
rect 514 193 516 208
rect 524 207 533 209
rect 524 204 526 207
rect 479 186 485 188
rect 479 184 481 186
rect 483 184 485 186
rect 479 182 485 184
rect 480 179 482 182
rect 406 165 408 170
rect 416 165 418 170
rect 423 165 425 170
rect 359 160 378 162
rect 433 162 435 170
rect 440 166 442 170
rect 450 162 452 172
rect 490 178 492 192
rect 497 191 509 193
rect 497 185 503 187
rect 497 183 499 185
rect 501 183 503 185
rect 497 181 503 183
rect 497 178 499 181
rect 507 178 509 191
rect 514 191 520 193
rect 514 189 516 191
rect 518 189 520 191
rect 514 187 520 189
rect 514 178 516 187
rect 524 178 526 196
rect 480 165 482 170
rect 490 165 492 170
rect 497 165 499 170
rect 433 160 452 162
rect 507 162 509 170
rect 514 166 516 170
rect 524 162 526 172
rect 507 160 526 162
rect -22 141 -20 146
rect -12 138 -10 143
rect -2 138 0 143
rect 18 143 20 147
rect 31 145 33 150
rect 38 145 40 150
rect 61 154 86 156
rect 61 146 63 154
rect 74 146 76 150
rect 84 146 86 154
rect 94 149 96 154
rect 101 149 103 154
rect 58 144 63 146
rect 58 141 60 144
rect -22 129 -20 132
rect -12 129 -10 132
rect -22 127 -16 129
rect -22 125 -20 127
rect -18 125 -16 127
rect -22 123 -16 125
rect -12 127 -6 129
rect -12 125 -10 127
rect -8 125 -6 127
rect -12 123 -6 125
rect -22 120 -20 123
rect -9 113 -7 123
rect -2 122 0 132
rect 18 129 20 134
rect 31 129 33 134
rect 18 127 24 129
rect 18 125 20 127
rect 22 125 24 127
rect 18 123 24 125
rect 28 127 34 129
rect 28 125 30 127
rect 32 125 34 127
rect 28 123 34 125
rect -2 120 4 122
rect -2 118 0 120
rect 2 118 4 120
rect 18 119 20 123
rect -2 116 4 118
rect -2 113 0 116
rect -22 97 -20 102
rect 28 112 30 123
rect 38 121 40 134
rect 122 143 124 147
rect 135 145 137 150
rect 142 145 144 150
rect 165 154 190 156
rect 165 146 167 154
rect 178 146 180 150
rect 188 146 190 154
rect 198 149 200 154
rect 205 149 207 154
rect 74 134 76 137
rect 67 132 76 134
rect 84 133 86 137
rect 94 134 96 137
rect 58 124 60 132
rect 67 130 69 132
rect 71 130 76 132
rect 67 128 76 130
rect 92 132 96 134
rect 92 129 94 132
rect 74 124 76 128
rect 88 127 94 129
rect 101 128 103 137
rect 162 144 167 146
rect 162 141 164 144
rect 122 129 124 134
rect 135 129 137 134
rect 88 125 90 127
rect 92 125 94 127
rect 55 122 68 124
rect 74 122 84 124
rect 88 123 94 125
rect 55 121 57 122
rect 38 119 44 121
rect 38 117 40 119
rect 42 117 44 119
rect 38 115 44 117
rect 51 119 57 121
rect 66 119 68 122
rect 82 119 84 122
rect 92 119 94 123
rect 98 126 104 128
rect 98 124 100 126
rect 102 124 104 126
rect 98 122 104 124
rect 102 119 104 122
rect 122 127 128 129
rect 122 125 124 127
rect 126 125 128 127
rect 122 123 128 125
rect 132 127 138 129
rect 132 125 134 127
rect 136 125 138 127
rect 132 123 138 125
rect 122 119 124 123
rect 51 117 53 119
rect 55 117 57 119
rect 51 115 57 117
rect 38 112 40 115
rect 18 97 20 101
rect 28 94 30 99
rect 38 94 40 99
rect -9 88 -7 92
rect -2 88 0 92
rect 82 97 84 101
rect 92 97 94 101
rect 66 88 68 92
rect 132 112 134 123
rect 142 121 144 134
rect 235 145 237 150
rect 242 145 244 150
rect 359 154 378 156
rect 178 134 180 137
rect 171 132 180 134
rect 188 133 190 137
rect 198 134 200 137
rect 162 124 164 132
rect 171 130 173 132
rect 175 130 180 132
rect 171 128 180 130
rect 196 132 200 134
rect 196 129 198 132
rect 178 124 180 128
rect 192 127 198 129
rect 205 128 207 137
rect 255 143 257 147
rect 332 146 334 151
rect 342 146 344 151
rect 349 146 351 151
rect 359 146 361 154
rect 366 146 368 150
rect 283 138 285 143
rect 293 138 295 143
rect 303 141 305 146
rect 192 125 194 127
rect 196 125 198 127
rect 159 122 172 124
rect 178 122 188 124
rect 192 123 198 125
rect 159 121 161 122
rect 142 119 148 121
rect 142 117 144 119
rect 146 117 148 119
rect 142 115 148 117
rect 155 119 161 121
rect 170 119 172 122
rect 186 119 188 122
rect 196 119 198 123
rect 202 126 208 128
rect 202 124 204 126
rect 206 124 208 126
rect 202 122 208 124
rect 206 119 208 122
rect 235 121 237 134
rect 242 129 244 134
rect 255 129 257 134
rect 376 144 378 154
rect 433 154 452 156
rect 406 146 408 151
rect 416 146 418 151
rect 423 146 425 151
rect 433 146 435 154
rect 440 146 442 150
rect 332 134 334 137
rect 331 132 337 134
rect 241 127 247 129
rect 241 125 243 127
rect 245 125 247 127
rect 241 123 247 125
rect 251 127 257 129
rect 251 125 253 127
rect 255 125 257 127
rect 251 123 257 125
rect 231 119 237 121
rect 155 117 157 119
rect 159 117 161 119
rect 155 115 161 117
rect 142 112 144 115
rect 122 97 124 101
rect 132 94 134 99
rect 142 94 144 99
rect 102 88 104 92
rect 186 97 188 101
rect 196 97 198 101
rect 170 88 172 92
rect 231 117 233 119
rect 235 117 237 119
rect 231 115 237 117
rect 235 112 237 115
rect 245 112 247 123
rect 255 119 257 123
rect 283 122 285 132
rect 293 129 295 132
rect 303 129 305 132
rect 289 127 295 129
rect 289 125 291 127
rect 293 125 295 127
rect 289 123 295 125
rect 299 127 305 129
rect 331 130 333 132
rect 335 130 337 132
rect 331 128 337 130
rect 299 125 301 127
rect 303 125 305 127
rect 299 123 305 125
rect 279 120 285 122
rect 279 118 281 120
rect 283 118 285 120
rect 279 116 285 118
rect 283 113 285 116
rect 290 113 292 123
rect 303 120 305 123
rect 235 94 237 99
rect 245 94 247 99
rect 255 97 257 101
rect 206 88 208 92
rect 332 110 334 128
rect 342 124 344 138
rect 349 135 351 138
rect 349 133 355 135
rect 349 131 351 133
rect 353 131 355 133
rect 349 129 355 131
rect 359 125 361 138
rect 339 122 345 124
rect 339 120 341 122
rect 343 120 345 122
rect 339 118 345 120
rect 349 123 361 125
rect 366 134 368 138
rect 366 132 372 134
rect 366 130 368 132
rect 370 130 372 132
rect 366 123 372 130
rect 303 97 305 102
rect 283 88 285 92
rect 290 88 292 92
rect 342 108 344 118
rect 349 108 351 123
rect 356 117 362 119
rect 356 115 358 117
rect 360 115 362 117
rect 356 113 362 115
rect 359 108 361 113
rect 366 108 368 123
rect 376 120 378 138
rect 450 144 452 154
rect 507 154 526 156
rect 480 146 482 151
rect 490 146 492 151
rect 497 146 499 151
rect 507 146 509 154
rect 514 146 516 150
rect 406 134 408 137
rect 405 132 411 134
rect 405 130 407 132
rect 409 130 411 132
rect 405 128 411 130
rect 376 109 378 112
rect 406 110 408 128
rect 416 124 418 138
rect 423 135 425 138
rect 423 133 429 135
rect 423 131 425 133
rect 427 131 429 133
rect 423 129 429 131
rect 433 125 435 138
rect 413 122 419 124
rect 413 120 415 122
rect 417 120 419 122
rect 413 118 419 120
rect 423 123 435 125
rect 440 129 442 138
rect 440 127 446 129
rect 440 125 442 127
rect 444 125 446 127
rect 440 123 446 125
rect 376 107 385 109
rect 379 105 381 107
rect 383 105 385 107
rect 379 103 385 105
rect 416 108 418 118
rect 423 108 425 123
rect 430 117 436 119
rect 430 115 432 117
rect 434 115 436 117
rect 430 113 436 115
rect 433 108 435 113
rect 440 108 442 123
rect 450 120 452 138
rect 524 144 526 154
rect 480 134 482 137
rect 479 132 485 134
rect 479 130 481 132
rect 483 130 485 132
rect 479 128 485 130
rect 450 109 452 112
rect 480 110 482 128
rect 490 124 492 138
rect 497 135 499 138
rect 497 133 503 135
rect 497 131 499 133
rect 501 131 503 133
rect 497 129 503 131
rect 507 125 509 138
rect 487 122 493 124
rect 487 120 489 122
rect 491 120 493 122
rect 487 118 493 120
rect 497 123 509 125
rect 514 129 516 138
rect 514 127 520 129
rect 514 125 516 127
rect 518 125 520 127
rect 514 123 520 125
rect 450 107 459 109
rect 453 105 455 107
rect 457 105 459 107
rect 453 103 459 105
rect 490 108 492 118
rect 497 108 499 123
rect 504 117 510 119
rect 504 115 506 117
rect 508 115 510 117
rect 504 113 510 115
rect 507 108 509 113
rect 514 108 516 123
rect 524 120 526 138
rect 524 109 526 112
rect 524 107 533 109
rect 527 105 529 107
rect 531 105 533 107
rect 527 103 533 105
rect 332 88 334 92
rect 342 88 344 92
rect 349 88 351 92
rect 359 88 361 92
rect 366 88 368 92
rect 406 88 408 92
rect 416 88 418 92
rect 423 88 425 92
rect 433 88 435 92
rect 440 88 442 92
rect 480 88 482 92
rect 490 88 492 92
rect 497 88 499 92
rect 507 88 509 92
rect 514 88 516 92
rect -9 80 -7 84
rect -2 80 0 84
rect -22 70 -20 75
rect 66 80 68 84
rect 18 71 20 75
rect 28 73 30 78
rect 38 73 40 78
rect -22 49 -20 52
rect -9 49 -7 59
rect -2 56 0 59
rect -2 54 4 56
rect -2 52 0 54
rect 2 52 4 54
rect -2 50 4 52
rect -22 47 -16 49
rect -22 45 -20 47
rect -18 45 -16 47
rect -22 43 -16 45
rect -12 47 -6 49
rect -12 45 -10 47
rect -8 45 -6 47
rect -12 43 -6 45
rect -22 40 -20 43
rect -12 40 -10 43
rect -2 40 0 50
rect 18 49 20 53
rect 28 49 30 60
rect 38 57 40 60
rect 38 55 44 57
rect 38 53 40 55
rect 42 53 44 55
rect 38 51 44 53
rect 51 55 57 57
rect 51 53 53 55
rect 55 53 57 55
rect 102 80 104 84
rect 82 71 84 75
rect 92 71 94 75
rect 170 80 172 84
rect 122 71 124 75
rect 132 73 134 78
rect 142 73 144 78
rect 51 51 57 53
rect 18 47 24 49
rect 18 45 20 47
rect 22 45 24 47
rect 18 43 24 45
rect 28 47 34 49
rect 28 45 30 47
rect 32 45 34 47
rect 28 43 34 45
rect 18 38 20 43
rect 31 38 33 43
rect 38 38 40 51
rect 55 50 57 51
rect 66 50 68 53
rect 82 50 84 53
rect 55 48 68 50
rect 74 48 84 50
rect 92 49 94 53
rect 102 50 104 53
rect 58 40 60 48
rect 74 44 76 48
rect 67 42 76 44
rect 88 47 94 49
rect 88 45 90 47
rect 92 45 94 47
rect 88 43 94 45
rect 98 48 104 50
rect 98 46 100 48
rect 102 46 104 48
rect 98 44 104 46
rect 122 49 124 53
rect 132 49 134 60
rect 142 57 144 60
rect 142 55 148 57
rect 142 53 144 55
rect 146 53 148 55
rect 142 51 148 53
rect 155 55 161 57
rect 155 53 157 55
rect 159 53 161 55
rect 206 80 208 84
rect 186 71 188 75
rect 196 71 198 75
rect 283 80 285 84
rect 290 80 292 84
rect 235 73 237 78
rect 245 73 247 78
rect 255 71 257 75
rect 235 57 237 60
rect 231 55 237 57
rect 231 53 233 55
rect 235 53 237 55
rect 155 51 161 53
rect 122 47 128 49
rect 122 45 124 47
rect 126 45 128 47
rect 67 40 69 42
rect 71 40 76 42
rect -22 26 -20 31
rect -12 29 -10 34
rect -2 29 0 34
rect 18 25 20 29
rect 67 38 76 40
rect 92 40 94 43
rect 74 35 76 38
rect 84 35 86 39
rect 92 38 96 40
rect 94 35 96 38
rect 101 35 103 44
rect 122 43 128 45
rect 132 47 138 49
rect 132 45 134 47
rect 136 45 138 47
rect 132 43 138 45
rect 122 38 124 43
rect 135 38 137 43
rect 142 38 144 51
rect 159 50 161 51
rect 170 50 172 53
rect 186 50 188 53
rect 159 48 172 50
rect 178 48 188 50
rect 196 49 198 53
rect 206 50 208 53
rect 231 51 237 53
rect 162 40 164 48
rect 178 44 180 48
rect 171 42 180 44
rect 192 47 198 49
rect 192 45 194 47
rect 196 45 198 47
rect 192 43 198 45
rect 202 48 208 50
rect 202 46 204 48
rect 206 46 208 48
rect 202 44 208 46
rect 171 40 173 42
rect 175 40 180 42
rect 58 28 60 31
rect 31 22 33 27
rect 38 22 40 27
rect 58 26 63 28
rect 61 18 63 26
rect 74 22 76 26
rect 84 18 86 26
rect 122 25 124 29
rect 171 38 180 40
rect 196 40 198 43
rect 178 35 180 38
rect 188 35 190 39
rect 196 38 200 40
rect 198 35 200 38
rect 205 35 207 44
rect 235 38 237 51
rect 245 49 247 60
rect 332 80 334 84
rect 342 80 344 84
rect 349 80 351 84
rect 359 80 361 84
rect 366 80 368 84
rect 406 80 408 84
rect 416 80 418 84
rect 423 80 425 84
rect 433 80 435 84
rect 440 80 442 84
rect 480 80 482 84
rect 490 80 492 84
rect 497 80 499 84
rect 507 80 509 84
rect 514 80 516 84
rect 303 70 305 75
rect 283 56 285 59
rect 279 54 285 56
rect 255 49 257 53
rect 279 52 281 54
rect 283 52 285 54
rect 279 50 285 52
rect 241 47 247 49
rect 241 45 243 47
rect 245 45 247 47
rect 241 43 247 45
rect 251 47 257 49
rect 251 45 253 47
rect 255 45 257 47
rect 251 43 257 45
rect 242 38 244 43
rect 255 38 257 43
rect 283 40 285 50
rect 290 49 292 59
rect 379 67 385 69
rect 379 65 381 67
rect 383 65 385 67
rect 303 49 305 52
rect 289 47 295 49
rect 289 45 291 47
rect 293 45 295 47
rect 289 43 295 45
rect 299 47 305 49
rect 299 45 301 47
rect 303 45 305 47
rect 299 43 305 45
rect 332 44 334 62
rect 342 54 344 64
rect 339 52 345 54
rect 339 50 341 52
rect 343 50 345 52
rect 339 48 345 50
rect 349 49 351 64
rect 359 59 361 64
rect 356 57 362 59
rect 356 55 358 57
rect 360 55 362 57
rect 356 53 362 55
rect 366 49 368 64
rect 376 63 385 65
rect 376 60 378 63
rect 453 67 459 69
rect 453 65 455 67
rect 457 65 459 67
rect 293 40 295 43
rect 303 40 305 43
rect 331 42 337 44
rect 331 40 333 42
rect 335 40 337 42
rect 162 28 164 31
rect 94 18 96 23
rect 101 18 103 23
rect 61 16 86 18
rect 135 22 137 27
rect 142 22 144 27
rect 162 26 167 28
rect 165 18 167 26
rect 178 22 180 26
rect 188 18 190 26
rect 198 18 200 23
rect 205 18 207 23
rect 235 22 237 27
rect 242 22 244 27
rect 165 16 190 18
rect 255 25 257 29
rect 283 29 285 34
rect 293 29 295 34
rect 331 38 337 40
rect 332 35 334 38
rect 303 26 305 31
rect 342 34 344 48
rect 349 47 361 49
rect 349 41 355 43
rect 349 39 351 41
rect 353 39 355 41
rect 349 37 355 39
rect 349 34 351 37
rect 359 34 361 47
rect 366 42 372 49
rect 366 40 368 42
rect 370 40 372 42
rect 366 38 372 40
rect 366 34 368 38
rect 376 34 378 52
rect 406 44 408 62
rect 416 54 418 64
rect 413 52 419 54
rect 413 50 415 52
rect 417 50 419 52
rect 413 48 419 50
rect 423 49 425 64
rect 433 59 435 64
rect 430 57 436 59
rect 430 55 432 57
rect 434 55 436 57
rect 430 53 436 55
rect 440 49 442 64
rect 450 63 459 65
rect 450 60 452 63
rect 527 67 533 69
rect 527 65 529 67
rect 531 65 533 67
rect 405 42 411 44
rect 405 40 407 42
rect 409 40 411 42
rect 405 38 411 40
rect 406 35 408 38
rect 332 21 334 26
rect 342 21 344 26
rect 349 21 351 26
rect 359 18 361 26
rect 366 22 368 26
rect 376 18 378 28
rect 416 34 418 48
rect 423 47 435 49
rect 423 41 429 43
rect 423 39 425 41
rect 427 39 429 41
rect 423 37 429 39
rect 423 34 425 37
rect 433 34 435 47
rect 440 47 446 49
rect 440 45 442 47
rect 444 45 446 47
rect 440 43 446 45
rect 440 34 442 43
rect 450 34 452 52
rect 480 44 482 62
rect 490 54 492 64
rect 487 52 493 54
rect 487 50 489 52
rect 491 50 493 52
rect 487 48 493 50
rect 497 49 499 64
rect 507 59 509 64
rect 504 57 510 59
rect 504 55 506 57
rect 508 55 510 57
rect 504 53 510 55
rect 514 49 516 64
rect 524 63 533 65
rect 524 60 526 63
rect 479 42 485 44
rect 479 40 481 42
rect 483 40 485 42
rect 479 38 485 40
rect 480 35 482 38
rect 406 21 408 26
rect 416 21 418 26
rect 423 21 425 26
rect 359 16 378 18
rect 433 18 435 26
rect 440 22 442 26
rect 450 18 452 28
rect 490 34 492 48
rect 497 47 509 49
rect 497 41 503 43
rect 497 39 499 41
rect 501 39 503 41
rect 497 37 503 39
rect 497 34 499 37
rect 507 34 509 47
rect 514 47 520 49
rect 514 45 516 47
rect 518 45 520 47
rect 514 43 520 45
rect 514 34 516 43
rect 524 34 526 52
rect 480 21 482 26
rect 490 21 492 26
rect 497 21 499 26
rect 433 16 452 18
rect 507 18 509 26
rect 514 22 516 26
rect 524 18 526 28
rect 507 16 526 18
<< ndif >>
rect -18 293 -12 295
rect -18 291 -16 293
rect -14 291 -12 293
rect -18 289 -12 291
rect 1 293 7 295
rect 22 297 29 299
rect 22 295 24 297
rect 26 295 29 297
rect 1 291 3 293
rect 5 291 7 293
rect 1 289 7 291
rect -18 285 -14 289
rect -27 282 -22 285
rect -29 280 -22 282
rect -29 278 -27 280
rect -25 278 -22 280
rect -29 276 -22 278
rect -20 282 -14 285
rect 2 282 7 289
rect 22 289 29 295
rect 105 297 111 299
rect 105 295 107 297
rect 109 295 111 297
rect 105 293 111 295
rect 126 297 133 299
rect 126 295 128 297
rect 130 295 133 297
rect 89 290 94 293
rect 22 287 31 289
rect -20 276 -12 282
rect -10 280 -2 282
rect -10 278 -7 280
rect -5 278 -2 280
rect -10 276 -2 278
rect 0 276 7 282
rect 11 285 18 287
rect 11 283 13 285
rect 15 283 18 285
rect 11 281 18 283
rect 13 278 18 281
rect 20 278 31 287
rect 33 278 38 289
rect 40 287 47 289
rect 40 285 43 287
rect 45 285 47 287
rect 65 288 74 290
rect 65 286 67 288
rect 69 286 74 288
rect 65 285 74 286
rect 40 283 47 285
rect 40 278 45 283
rect 53 282 58 285
rect 51 280 58 282
rect 51 278 53 280
rect 55 278 58 280
rect 51 276 58 278
rect 60 281 74 285
rect 76 285 84 290
rect 76 283 79 285
rect 81 283 84 285
rect 76 281 84 283
rect 86 287 94 290
rect 86 285 89 287
rect 91 285 94 287
rect 86 281 94 285
rect 96 281 101 293
rect 103 281 111 293
rect 126 289 133 295
rect 209 297 215 299
rect 209 295 211 297
rect 213 295 215 297
rect 209 293 215 295
rect 246 297 253 299
rect 246 295 249 297
rect 251 295 253 297
rect 193 290 198 293
rect 126 287 135 289
rect 115 285 122 287
rect 115 283 117 285
rect 119 283 122 285
rect 115 281 122 283
rect 60 276 65 281
rect 117 278 122 281
rect 124 278 135 287
rect 137 278 142 289
rect 144 287 151 289
rect 144 285 147 287
rect 149 285 151 287
rect 169 288 178 290
rect 169 286 171 288
rect 173 286 178 288
rect 169 285 178 286
rect 144 283 151 285
rect 144 278 149 283
rect 157 282 162 285
rect 155 280 162 282
rect 155 278 157 280
rect 159 278 162 280
rect 155 276 162 278
rect 164 281 178 285
rect 180 285 188 290
rect 180 283 183 285
rect 185 283 188 285
rect 180 281 188 283
rect 190 287 198 290
rect 190 285 193 287
rect 195 285 198 287
rect 190 281 198 285
rect 200 281 205 293
rect 207 281 215 293
rect 246 289 253 295
rect 276 293 282 295
rect 276 291 278 293
rect 280 291 282 293
rect 228 287 235 289
rect 228 285 230 287
rect 232 285 235 287
rect 228 283 235 285
rect 164 276 169 281
rect 230 278 235 283
rect 237 278 242 289
rect 244 287 253 289
rect 276 289 282 291
rect 295 293 301 295
rect 295 291 297 293
rect 299 291 301 293
rect 295 289 301 291
rect 244 278 255 287
rect 257 285 264 287
rect 257 283 260 285
rect 262 283 264 285
rect 257 281 264 283
rect 276 282 281 289
rect 297 285 301 289
rect 327 287 332 290
rect 325 285 332 287
rect 297 282 303 285
rect 257 278 262 281
rect 276 276 283 282
rect 285 280 293 282
rect 285 278 288 280
rect 290 278 293 280
rect 285 276 293 278
rect 295 276 303 282
rect 305 282 310 285
rect 325 283 327 285
rect 329 283 332 285
rect 305 280 312 282
rect 325 281 332 283
rect 334 288 342 290
rect 334 286 337 288
rect 339 286 342 288
rect 334 282 342 286
rect 344 282 349 290
rect 351 288 359 290
rect 351 286 354 288
rect 356 286 359 288
rect 351 282 359 286
rect 361 282 366 290
rect 368 288 374 290
rect 368 286 376 288
rect 368 284 371 286
rect 373 284 376 286
rect 368 282 376 284
rect 378 286 385 288
rect 401 287 406 290
rect 378 284 381 286
rect 383 284 385 286
rect 378 282 385 284
rect 399 285 406 287
rect 399 283 401 285
rect 403 283 406 285
rect 334 281 339 282
rect 305 278 308 280
rect 310 278 312 280
rect 305 276 312 278
rect 399 281 406 283
rect 408 288 416 290
rect 408 286 411 288
rect 413 286 416 288
rect 408 282 416 286
rect 418 282 423 290
rect 425 288 433 290
rect 425 286 428 288
rect 430 286 433 288
rect 425 282 433 286
rect 435 282 440 290
rect 442 288 448 290
rect 442 286 450 288
rect 442 284 445 286
rect 447 284 450 286
rect 442 282 450 284
rect 452 286 459 288
rect 475 287 480 290
rect 452 284 455 286
rect 457 284 459 286
rect 452 282 459 284
rect 473 285 480 287
rect 473 283 475 285
rect 477 283 480 285
rect 408 281 413 282
rect 473 281 480 283
rect 482 288 490 290
rect 482 286 485 288
rect 487 286 490 288
rect 482 282 490 286
rect 492 282 497 290
rect 499 288 507 290
rect 499 286 502 288
rect 504 286 507 288
rect 499 282 507 286
rect 509 282 514 290
rect 516 288 522 290
rect 516 286 524 288
rect 516 284 519 286
rect 521 284 524 286
rect 516 282 524 284
rect 526 286 533 288
rect 526 284 529 286
rect 531 284 533 286
rect 526 282 533 284
rect 482 281 487 282
rect -29 182 -22 184
rect -29 180 -27 182
rect -25 180 -22 182
rect -29 178 -22 180
rect -27 175 -22 178
rect -20 178 -12 184
rect -10 182 -2 184
rect -10 180 -7 182
rect -5 180 -2 182
rect -10 178 -2 180
rect 0 178 7 184
rect 51 182 58 184
rect 13 179 18 182
rect -20 175 -14 178
rect -18 171 -14 175
rect 2 171 7 178
rect 11 177 18 179
rect 11 175 13 177
rect 15 175 18 177
rect 11 173 18 175
rect 20 173 31 182
rect -18 169 -12 171
rect -18 167 -16 169
rect -14 167 -12 169
rect -18 165 -12 167
rect 1 169 7 171
rect 22 171 31 173
rect 33 171 38 182
rect 40 177 45 182
rect 51 180 53 182
rect 55 180 58 182
rect 51 178 58 180
rect 40 175 47 177
rect 53 175 58 178
rect 60 179 65 184
rect 155 182 162 184
rect 117 179 122 182
rect 60 175 74 179
rect 40 173 43 175
rect 45 173 47 175
rect 40 171 47 173
rect 65 174 74 175
rect 65 172 67 174
rect 69 172 74 174
rect 1 167 3 169
rect 5 167 7 169
rect 1 165 7 167
rect 22 165 29 171
rect 65 170 74 172
rect 76 177 84 179
rect 76 175 79 177
rect 81 175 84 177
rect 76 170 84 175
rect 86 175 94 179
rect 86 173 89 175
rect 91 173 94 175
rect 86 170 94 173
rect 22 163 24 165
rect 26 163 29 165
rect 22 161 29 163
rect 89 167 94 170
rect 96 167 101 179
rect 103 167 111 179
rect 115 177 122 179
rect 115 175 117 177
rect 119 175 122 177
rect 115 173 122 175
rect 124 173 135 182
rect 126 171 135 173
rect 137 171 142 182
rect 144 177 149 182
rect 155 180 157 182
rect 159 180 162 182
rect 155 178 162 180
rect 144 175 151 177
rect 157 175 162 178
rect 164 179 169 184
rect 164 175 178 179
rect 144 173 147 175
rect 149 173 151 175
rect 144 171 151 173
rect 169 174 178 175
rect 169 172 171 174
rect 173 172 178 174
rect 105 165 111 167
rect 105 163 107 165
rect 109 163 111 165
rect 105 161 111 163
rect 126 165 133 171
rect 169 170 178 172
rect 180 177 188 179
rect 180 175 183 177
rect 185 175 188 177
rect 180 170 188 175
rect 190 175 198 179
rect 190 173 193 175
rect 195 173 198 175
rect 190 170 198 173
rect 126 163 128 165
rect 130 163 133 165
rect 126 161 133 163
rect 193 167 198 170
rect 200 167 205 179
rect 207 167 215 179
rect 230 177 235 182
rect 228 175 235 177
rect 228 173 230 175
rect 232 173 235 175
rect 228 171 235 173
rect 237 171 242 182
rect 244 173 255 182
rect 257 179 262 182
rect 257 177 264 179
rect 257 175 260 177
rect 262 175 264 177
rect 257 173 264 175
rect 276 178 283 184
rect 285 182 293 184
rect 285 180 288 182
rect 290 180 293 182
rect 285 178 293 180
rect 295 178 303 184
rect 244 171 253 173
rect 209 165 215 167
rect 209 163 211 165
rect 213 163 215 165
rect 209 161 215 163
rect 246 165 253 171
rect 276 171 281 178
rect 297 175 303 178
rect 305 182 312 184
rect 305 180 308 182
rect 310 180 312 182
rect 305 178 312 180
rect 305 175 310 178
rect 325 177 332 179
rect 325 175 327 177
rect 329 175 332 177
rect 297 171 301 175
rect 276 169 282 171
rect 276 167 278 169
rect 280 167 282 169
rect 246 163 249 165
rect 251 163 253 165
rect 246 161 253 163
rect 276 165 282 167
rect 295 169 301 171
rect 325 173 332 175
rect 327 170 332 173
rect 334 178 339 179
rect 334 174 342 178
rect 334 172 337 174
rect 339 172 342 174
rect 334 170 342 172
rect 344 170 349 178
rect 351 174 359 178
rect 351 172 354 174
rect 356 172 359 174
rect 351 170 359 172
rect 361 170 366 178
rect 368 176 376 178
rect 368 174 371 176
rect 373 174 376 176
rect 368 172 376 174
rect 378 176 385 178
rect 378 174 381 176
rect 383 174 385 176
rect 378 172 385 174
rect 399 177 406 179
rect 399 175 401 177
rect 403 175 406 177
rect 399 173 406 175
rect 368 170 374 172
rect 295 167 297 169
rect 299 167 301 169
rect 295 165 301 167
rect 401 170 406 173
rect 408 178 413 179
rect 408 174 416 178
rect 408 172 411 174
rect 413 172 416 174
rect 408 170 416 172
rect 418 170 423 178
rect 425 174 433 178
rect 425 172 428 174
rect 430 172 433 174
rect 425 170 433 172
rect 435 170 440 178
rect 442 176 450 178
rect 442 174 445 176
rect 447 174 450 176
rect 442 172 450 174
rect 452 176 459 178
rect 452 174 455 176
rect 457 174 459 176
rect 452 172 459 174
rect 473 177 480 179
rect 473 175 475 177
rect 477 175 480 177
rect 473 173 480 175
rect 442 170 448 172
rect 475 170 480 173
rect 482 178 487 179
rect 482 174 490 178
rect 482 172 485 174
rect 487 172 490 174
rect 482 170 490 172
rect 492 170 497 178
rect 499 174 507 178
rect 499 172 502 174
rect 504 172 507 174
rect 499 170 507 172
rect 509 170 514 178
rect 516 176 524 178
rect 516 174 519 176
rect 521 174 524 176
rect 516 172 524 174
rect 526 176 533 178
rect 526 174 529 176
rect 531 174 533 176
rect 526 172 533 174
rect 516 170 522 172
rect -18 149 -12 151
rect -18 147 -16 149
rect -14 147 -12 149
rect -18 145 -12 147
rect 1 149 7 151
rect 22 153 29 155
rect 22 151 24 153
rect 26 151 29 153
rect 1 147 3 149
rect 5 147 7 149
rect 1 145 7 147
rect -18 141 -14 145
rect -27 138 -22 141
rect -29 136 -22 138
rect -29 134 -27 136
rect -25 134 -22 136
rect -29 132 -22 134
rect -20 138 -14 141
rect 2 138 7 145
rect 22 145 29 151
rect 105 153 111 155
rect 105 151 107 153
rect 109 151 111 153
rect 105 149 111 151
rect 126 153 133 155
rect 126 151 128 153
rect 130 151 133 153
rect 89 146 94 149
rect 22 143 31 145
rect -20 132 -12 138
rect -10 136 -2 138
rect -10 134 -7 136
rect -5 134 -2 136
rect -10 132 -2 134
rect 0 132 7 138
rect 11 141 18 143
rect 11 139 13 141
rect 15 139 18 141
rect 11 137 18 139
rect 13 134 18 137
rect 20 134 31 143
rect 33 134 38 145
rect 40 143 47 145
rect 40 141 43 143
rect 45 141 47 143
rect 65 144 74 146
rect 65 142 67 144
rect 69 142 74 144
rect 65 141 74 142
rect 40 139 47 141
rect 40 134 45 139
rect 53 138 58 141
rect 51 136 58 138
rect 51 134 53 136
rect 55 134 58 136
rect 51 132 58 134
rect 60 137 74 141
rect 76 141 84 146
rect 76 139 79 141
rect 81 139 84 141
rect 76 137 84 139
rect 86 143 94 146
rect 86 141 89 143
rect 91 141 94 143
rect 86 137 94 141
rect 96 137 101 149
rect 103 137 111 149
rect 126 145 133 151
rect 209 153 215 155
rect 209 151 211 153
rect 213 151 215 153
rect 209 149 215 151
rect 246 153 253 155
rect 246 151 249 153
rect 251 151 253 153
rect 193 146 198 149
rect 126 143 135 145
rect 115 141 122 143
rect 115 139 117 141
rect 119 139 122 141
rect 115 137 122 139
rect 60 132 65 137
rect 117 134 122 137
rect 124 134 135 143
rect 137 134 142 145
rect 144 143 151 145
rect 144 141 147 143
rect 149 141 151 143
rect 169 144 178 146
rect 169 142 171 144
rect 173 142 178 144
rect 169 141 178 142
rect 144 139 151 141
rect 144 134 149 139
rect 157 138 162 141
rect 155 136 162 138
rect 155 134 157 136
rect 159 134 162 136
rect 155 132 162 134
rect 164 137 178 141
rect 180 141 188 146
rect 180 139 183 141
rect 185 139 188 141
rect 180 137 188 139
rect 190 143 198 146
rect 190 141 193 143
rect 195 141 198 143
rect 190 137 198 141
rect 200 137 205 149
rect 207 137 215 149
rect 246 145 253 151
rect 276 149 282 151
rect 276 147 278 149
rect 280 147 282 149
rect 228 143 235 145
rect 228 141 230 143
rect 232 141 235 143
rect 228 139 235 141
rect 164 132 169 137
rect 230 134 235 139
rect 237 134 242 145
rect 244 143 253 145
rect 276 145 282 147
rect 295 149 301 151
rect 295 147 297 149
rect 299 147 301 149
rect 295 145 301 147
rect 244 134 255 143
rect 257 141 264 143
rect 257 139 260 141
rect 262 139 264 141
rect 257 137 264 139
rect 276 138 281 145
rect 297 141 301 145
rect 327 143 332 146
rect 325 141 332 143
rect 297 138 303 141
rect 257 134 262 137
rect 276 132 283 138
rect 285 136 293 138
rect 285 134 288 136
rect 290 134 293 136
rect 285 132 293 134
rect 295 132 303 138
rect 305 138 310 141
rect 325 139 327 141
rect 329 139 332 141
rect 305 136 312 138
rect 325 137 332 139
rect 334 144 342 146
rect 334 142 337 144
rect 339 142 342 144
rect 334 138 342 142
rect 344 138 349 146
rect 351 144 359 146
rect 351 142 354 144
rect 356 142 359 144
rect 351 138 359 142
rect 361 138 366 146
rect 368 144 374 146
rect 368 142 376 144
rect 368 140 371 142
rect 373 140 376 142
rect 368 138 376 140
rect 378 142 385 144
rect 401 143 406 146
rect 378 140 381 142
rect 383 140 385 142
rect 378 138 385 140
rect 399 141 406 143
rect 399 139 401 141
rect 403 139 406 141
rect 334 137 339 138
rect 305 134 308 136
rect 310 134 312 136
rect 305 132 312 134
rect 399 137 406 139
rect 408 144 416 146
rect 408 142 411 144
rect 413 142 416 144
rect 408 138 416 142
rect 418 138 423 146
rect 425 144 433 146
rect 425 142 428 144
rect 430 142 433 144
rect 425 138 433 142
rect 435 138 440 146
rect 442 144 448 146
rect 442 142 450 144
rect 442 140 445 142
rect 447 140 450 142
rect 442 138 450 140
rect 452 142 459 144
rect 475 143 480 146
rect 452 140 455 142
rect 457 140 459 142
rect 452 138 459 140
rect 473 141 480 143
rect 473 139 475 141
rect 477 139 480 141
rect 408 137 413 138
rect 473 137 480 139
rect 482 144 490 146
rect 482 142 485 144
rect 487 142 490 144
rect 482 138 490 142
rect 492 138 497 146
rect 499 144 507 146
rect 499 142 502 144
rect 504 142 507 144
rect 499 138 507 142
rect 509 138 514 146
rect 516 144 522 146
rect 516 142 524 144
rect 516 140 519 142
rect 521 140 524 142
rect 516 138 524 140
rect 526 142 533 144
rect 526 140 529 142
rect 531 140 533 142
rect 526 138 533 140
rect 482 137 487 138
rect -29 38 -22 40
rect -29 36 -27 38
rect -25 36 -22 38
rect -29 34 -22 36
rect -27 31 -22 34
rect -20 34 -12 40
rect -10 38 -2 40
rect -10 36 -7 38
rect -5 36 -2 38
rect -10 34 -2 36
rect 0 34 7 40
rect 51 38 58 40
rect 13 35 18 38
rect -20 31 -14 34
rect -18 27 -14 31
rect 2 27 7 34
rect 11 33 18 35
rect 11 31 13 33
rect 15 31 18 33
rect 11 29 18 31
rect 20 29 31 38
rect -18 25 -12 27
rect -18 23 -16 25
rect -14 23 -12 25
rect -18 21 -12 23
rect 1 25 7 27
rect 22 27 31 29
rect 33 27 38 38
rect 40 33 45 38
rect 51 36 53 38
rect 55 36 58 38
rect 51 34 58 36
rect 40 31 47 33
rect 53 31 58 34
rect 60 35 65 40
rect 155 38 162 40
rect 117 35 122 38
rect 60 31 74 35
rect 40 29 43 31
rect 45 29 47 31
rect 40 27 47 29
rect 65 30 74 31
rect 65 28 67 30
rect 69 28 74 30
rect 1 23 3 25
rect 5 23 7 25
rect 1 21 7 23
rect 22 21 29 27
rect 65 26 74 28
rect 76 33 84 35
rect 76 31 79 33
rect 81 31 84 33
rect 76 26 84 31
rect 86 31 94 35
rect 86 29 89 31
rect 91 29 94 31
rect 86 26 94 29
rect 22 19 24 21
rect 26 19 29 21
rect 22 17 29 19
rect 89 23 94 26
rect 96 23 101 35
rect 103 23 111 35
rect 115 33 122 35
rect 115 31 117 33
rect 119 31 122 33
rect 115 29 122 31
rect 124 29 135 38
rect 126 27 135 29
rect 137 27 142 38
rect 144 33 149 38
rect 155 36 157 38
rect 159 36 162 38
rect 155 34 162 36
rect 144 31 151 33
rect 157 31 162 34
rect 164 35 169 40
rect 164 31 178 35
rect 144 29 147 31
rect 149 29 151 31
rect 144 27 151 29
rect 169 30 178 31
rect 169 28 171 30
rect 173 28 178 30
rect 105 21 111 23
rect 105 19 107 21
rect 109 19 111 21
rect 105 17 111 19
rect 126 21 133 27
rect 169 26 178 28
rect 180 33 188 35
rect 180 31 183 33
rect 185 31 188 33
rect 180 26 188 31
rect 190 31 198 35
rect 190 29 193 31
rect 195 29 198 31
rect 190 26 198 29
rect 126 19 128 21
rect 130 19 133 21
rect 126 17 133 19
rect 193 23 198 26
rect 200 23 205 35
rect 207 23 215 35
rect 230 33 235 38
rect 228 31 235 33
rect 228 29 230 31
rect 232 29 235 31
rect 228 27 235 29
rect 237 27 242 38
rect 244 29 255 38
rect 257 35 262 38
rect 257 33 264 35
rect 257 31 260 33
rect 262 31 264 33
rect 257 29 264 31
rect 276 34 283 40
rect 285 38 293 40
rect 285 36 288 38
rect 290 36 293 38
rect 285 34 293 36
rect 295 34 303 40
rect 244 27 253 29
rect 209 21 215 23
rect 209 19 211 21
rect 213 19 215 21
rect 209 17 215 19
rect 246 21 253 27
rect 276 27 281 34
rect 297 31 303 34
rect 305 38 312 40
rect 305 36 308 38
rect 310 36 312 38
rect 305 34 312 36
rect 305 31 310 34
rect 325 33 332 35
rect 325 31 327 33
rect 329 31 332 33
rect 297 27 301 31
rect 276 25 282 27
rect 276 23 278 25
rect 280 23 282 25
rect 246 19 249 21
rect 251 19 253 21
rect 246 17 253 19
rect 276 21 282 23
rect 295 25 301 27
rect 325 29 332 31
rect 327 26 332 29
rect 334 34 339 35
rect 334 30 342 34
rect 334 28 337 30
rect 339 28 342 30
rect 334 26 342 28
rect 344 26 349 34
rect 351 30 359 34
rect 351 28 354 30
rect 356 28 359 30
rect 351 26 359 28
rect 361 26 366 34
rect 368 32 376 34
rect 368 30 371 32
rect 373 30 376 32
rect 368 28 376 30
rect 378 32 385 34
rect 378 30 381 32
rect 383 30 385 32
rect 378 28 385 30
rect 399 33 406 35
rect 399 31 401 33
rect 403 31 406 33
rect 399 29 406 31
rect 368 26 374 28
rect 295 23 297 25
rect 299 23 301 25
rect 295 21 301 23
rect 401 26 406 29
rect 408 34 413 35
rect 408 30 416 34
rect 408 28 411 30
rect 413 28 416 30
rect 408 26 416 28
rect 418 26 423 34
rect 425 30 433 34
rect 425 28 428 30
rect 430 28 433 30
rect 425 26 433 28
rect 435 26 440 34
rect 442 32 450 34
rect 442 30 445 32
rect 447 30 450 32
rect 442 28 450 30
rect 452 32 459 34
rect 452 30 455 32
rect 457 30 459 32
rect 452 28 459 30
rect 473 33 480 35
rect 473 31 475 33
rect 477 31 480 33
rect 473 29 480 31
rect 442 26 448 28
rect 475 26 480 29
rect 482 34 487 35
rect 482 30 490 34
rect 482 28 485 30
rect 487 28 490 30
rect 482 26 490 28
rect 492 26 497 34
rect 499 30 507 34
rect 499 28 502 30
rect 504 28 507 30
rect 499 26 507 28
rect 509 26 514 34
rect 516 32 524 34
rect 516 30 519 32
rect 521 30 524 32
rect 516 28 524 30
rect 526 32 533 34
rect 526 30 529 32
rect 531 30 533 32
rect 526 28 533 30
rect 516 26 522 28
<< pdif >>
rect -27 259 -22 264
rect -29 257 -22 259
rect -29 255 -27 257
rect -25 255 -22 257
rect -29 250 -22 255
rect -29 248 -27 250
rect -25 248 -22 250
rect -29 246 -22 248
rect -20 257 -12 264
rect 11 261 18 263
rect 11 259 13 261
rect 15 259 18 261
rect -20 246 -9 257
rect -18 240 -9 246
rect -18 238 -16 240
rect -14 238 -9 240
rect -18 236 -9 238
rect -7 236 -2 257
rect 0 249 5 257
rect 11 254 18 259
rect 11 252 13 254
rect 15 252 18 254
rect 11 250 18 252
rect 0 247 7 249
rect 0 245 3 247
rect 5 245 7 247
rect 13 245 18 250
rect 20 256 26 263
rect 59 261 66 263
rect 59 259 61 261
rect 63 259 66 261
rect 59 257 66 259
rect 20 249 28 256
rect 20 247 23 249
rect 25 247 28 249
rect 20 245 28 247
rect 0 243 7 245
rect 0 236 5 243
rect 22 243 28 245
rect 30 254 38 256
rect 30 252 33 254
rect 35 252 38 254
rect 30 247 38 252
rect 30 245 33 247
rect 35 245 38 247
rect 30 243 38 245
rect 40 247 47 256
rect 40 245 43 247
rect 45 245 47 247
rect 40 243 47 245
rect 61 236 66 257
rect 68 247 82 263
rect 68 245 71 247
rect 73 245 82 247
rect 84 261 92 263
rect 84 259 87 261
rect 89 259 92 261
rect 84 254 92 259
rect 84 252 87 254
rect 89 252 92 254
rect 84 245 92 252
rect 94 254 102 263
rect 94 252 97 254
rect 99 252 102 254
rect 94 245 102 252
rect 68 240 80 245
rect 68 238 71 240
rect 73 238 80 240
rect 68 236 80 238
rect 97 236 102 245
rect 104 248 109 263
rect 115 261 122 263
rect 115 259 117 261
rect 119 259 122 261
rect 115 254 122 259
rect 115 252 117 254
rect 119 252 122 254
rect 115 250 122 252
rect 104 246 111 248
rect 104 244 107 246
rect 109 244 111 246
rect 117 245 122 250
rect 124 256 130 263
rect 163 261 170 263
rect 163 259 165 261
rect 167 259 170 261
rect 163 257 170 259
rect 124 249 132 256
rect 124 247 127 249
rect 129 247 132 249
rect 124 245 132 247
rect 104 242 111 244
rect 104 236 109 242
rect 126 243 132 245
rect 134 254 142 256
rect 134 252 137 254
rect 139 252 142 254
rect 134 247 142 252
rect 134 245 137 247
rect 139 245 142 247
rect 134 243 142 245
rect 144 247 151 256
rect 144 245 147 247
rect 149 245 151 247
rect 144 243 151 245
rect 165 236 170 257
rect 172 247 186 263
rect 172 245 175 247
rect 177 245 186 247
rect 188 261 196 263
rect 188 259 191 261
rect 193 259 196 261
rect 188 254 196 259
rect 188 252 191 254
rect 193 252 196 254
rect 188 245 196 252
rect 198 254 206 263
rect 198 252 201 254
rect 203 252 206 254
rect 198 245 206 252
rect 172 240 184 245
rect 172 238 175 240
rect 177 238 184 240
rect 172 236 184 238
rect 201 236 206 245
rect 208 248 213 263
rect 249 256 255 263
rect 208 246 215 248
rect 208 244 211 246
rect 213 244 215 246
rect 208 242 215 244
rect 228 247 235 256
rect 228 245 230 247
rect 232 245 235 247
rect 228 243 235 245
rect 237 254 245 256
rect 237 252 240 254
rect 242 252 245 254
rect 237 247 245 252
rect 237 245 240 247
rect 242 245 245 247
rect 237 243 245 245
rect 247 249 255 256
rect 247 247 250 249
rect 252 247 255 249
rect 247 245 255 247
rect 257 261 264 263
rect 257 259 260 261
rect 262 259 264 261
rect 257 254 264 259
rect 295 257 303 264
rect 257 252 260 254
rect 262 252 264 254
rect 257 250 264 252
rect 257 245 262 250
rect 278 249 283 257
rect 276 247 283 249
rect 276 245 278 247
rect 280 245 283 247
rect 247 243 253 245
rect 208 236 213 242
rect 276 243 283 245
rect 278 236 283 243
rect 285 236 290 257
rect 292 246 303 257
rect 305 259 310 264
rect 305 257 312 259
rect 305 255 308 257
rect 310 255 312 257
rect 305 250 312 255
rect 305 248 308 250
rect 310 248 312 250
rect 327 249 332 254
rect 305 246 312 248
rect 325 247 332 249
rect 292 240 301 246
rect 325 245 327 247
rect 329 245 332 247
rect 325 243 332 245
rect 292 238 297 240
rect 299 238 301 240
rect 292 236 301 238
rect 327 236 332 243
rect 334 252 339 254
rect 370 256 376 264
rect 378 262 385 264
rect 378 260 381 262
rect 383 260 385 262
rect 378 258 385 260
rect 378 256 383 258
rect 370 252 374 256
rect 334 240 342 252
rect 334 238 337 240
rect 339 238 342 240
rect 334 236 342 238
rect 344 236 349 252
rect 351 250 359 252
rect 351 248 354 250
rect 356 248 359 250
rect 351 236 359 248
rect 361 236 366 252
rect 368 248 374 252
rect 401 249 406 254
rect 368 240 375 248
rect 399 247 406 249
rect 399 245 401 247
rect 403 245 406 247
rect 399 243 406 245
rect 368 238 371 240
rect 373 238 375 240
rect 368 236 375 238
rect 401 236 406 243
rect 408 252 413 254
rect 444 256 450 264
rect 452 262 459 264
rect 452 260 455 262
rect 457 260 459 262
rect 452 258 459 260
rect 452 256 457 258
rect 444 252 448 256
rect 408 240 416 252
rect 408 238 411 240
rect 413 238 416 240
rect 408 236 416 238
rect 418 236 423 252
rect 425 250 433 252
rect 425 248 428 250
rect 430 248 433 250
rect 425 236 433 248
rect 435 236 440 252
rect 442 248 448 252
rect 475 249 480 254
rect 442 240 449 248
rect 473 247 480 249
rect 473 245 475 247
rect 477 245 480 247
rect 473 243 480 245
rect 442 238 445 240
rect 447 238 449 240
rect 442 236 449 238
rect 475 236 480 243
rect 482 252 487 254
rect 518 256 524 264
rect 526 262 533 264
rect 526 260 529 262
rect 531 260 533 262
rect 526 258 533 260
rect 526 256 531 258
rect 518 252 522 256
rect 482 240 490 252
rect 482 238 485 240
rect 487 238 490 240
rect 482 236 490 238
rect 492 236 497 252
rect 499 250 507 252
rect 499 248 502 250
rect 504 248 507 250
rect 499 236 507 248
rect 509 236 514 252
rect 516 248 522 252
rect 516 240 523 248
rect 516 238 519 240
rect 521 238 523 240
rect 516 236 523 238
rect -18 222 -9 224
rect -18 220 -16 222
rect -14 220 -9 222
rect -18 214 -9 220
rect -29 212 -22 214
rect -29 210 -27 212
rect -25 210 -22 212
rect -29 205 -22 210
rect -29 203 -27 205
rect -25 203 -22 205
rect -29 201 -22 203
rect -27 196 -22 201
rect -20 203 -9 214
rect -7 203 -2 224
rect 0 217 5 224
rect 0 215 7 217
rect 22 215 28 217
rect 0 213 3 215
rect 5 213 7 215
rect 0 211 7 213
rect 0 203 5 211
rect 13 210 18 215
rect 11 208 18 210
rect 11 206 13 208
rect 15 206 18 208
rect -20 196 -12 203
rect 11 201 18 206
rect 11 199 13 201
rect 15 199 18 201
rect 11 197 18 199
rect 20 213 28 215
rect 20 211 23 213
rect 25 211 28 213
rect 20 204 28 211
rect 30 215 38 217
rect 30 213 33 215
rect 35 213 38 215
rect 30 208 38 213
rect 30 206 33 208
rect 35 206 38 208
rect 30 204 38 206
rect 40 215 47 217
rect 40 213 43 215
rect 45 213 47 215
rect 40 204 47 213
rect 20 197 26 204
rect 61 203 66 224
rect 59 201 66 203
rect 59 199 61 201
rect 63 199 66 201
rect 59 197 66 199
rect 68 222 80 224
rect 68 220 71 222
rect 73 220 80 222
rect 68 215 80 220
rect 97 215 102 224
rect 68 213 71 215
rect 73 213 82 215
rect 68 197 82 213
rect 84 208 92 215
rect 84 206 87 208
rect 89 206 92 208
rect 84 201 92 206
rect 84 199 87 201
rect 89 199 92 201
rect 84 197 92 199
rect 94 208 102 215
rect 94 206 97 208
rect 99 206 102 208
rect 94 197 102 206
rect 104 218 109 224
rect 104 216 111 218
rect 104 214 107 216
rect 109 214 111 216
rect 126 215 132 217
rect 104 212 111 214
rect 104 197 109 212
rect 117 210 122 215
rect 115 208 122 210
rect 115 206 117 208
rect 119 206 122 208
rect 115 201 122 206
rect 115 199 117 201
rect 119 199 122 201
rect 115 197 122 199
rect 124 213 132 215
rect 124 211 127 213
rect 129 211 132 213
rect 124 204 132 211
rect 134 215 142 217
rect 134 213 137 215
rect 139 213 142 215
rect 134 208 142 213
rect 134 206 137 208
rect 139 206 142 208
rect 134 204 142 206
rect 144 215 151 217
rect 144 213 147 215
rect 149 213 151 215
rect 144 204 151 213
rect 124 197 130 204
rect 165 203 170 224
rect 163 201 170 203
rect 163 199 165 201
rect 167 199 170 201
rect 163 197 170 199
rect 172 222 184 224
rect 172 220 175 222
rect 177 220 184 222
rect 172 215 184 220
rect 201 215 206 224
rect 172 213 175 215
rect 177 213 186 215
rect 172 197 186 213
rect 188 208 196 215
rect 188 206 191 208
rect 193 206 196 208
rect 188 201 196 206
rect 188 199 191 201
rect 193 199 196 201
rect 188 197 196 199
rect 198 208 206 215
rect 198 206 201 208
rect 203 206 206 208
rect 198 197 206 206
rect 208 218 213 224
rect 208 216 215 218
rect 208 214 211 216
rect 213 214 215 216
rect 208 212 215 214
rect 228 215 235 217
rect 228 213 230 215
rect 232 213 235 215
rect 208 197 213 212
rect 228 204 235 213
rect 237 215 245 217
rect 237 213 240 215
rect 242 213 245 215
rect 237 208 245 213
rect 237 206 240 208
rect 242 206 245 208
rect 237 204 245 206
rect 247 215 253 217
rect 278 217 283 224
rect 276 215 283 217
rect 247 213 255 215
rect 247 211 250 213
rect 252 211 255 213
rect 247 204 255 211
rect 249 197 255 204
rect 257 210 262 215
rect 276 213 278 215
rect 280 213 283 215
rect 276 211 283 213
rect 257 208 264 210
rect 257 206 260 208
rect 262 206 264 208
rect 257 201 264 206
rect 278 203 283 211
rect 285 203 290 224
rect 292 222 301 224
rect 292 220 297 222
rect 299 220 301 222
rect 292 214 301 220
rect 327 217 332 224
rect 325 215 332 217
rect 292 203 303 214
rect 257 199 260 201
rect 262 199 264 201
rect 257 197 264 199
rect 295 196 303 203
rect 305 212 312 214
rect 305 210 308 212
rect 310 210 312 212
rect 325 213 327 215
rect 329 213 332 215
rect 325 211 332 213
rect 305 205 312 210
rect 327 206 332 211
rect 334 222 342 224
rect 334 220 337 222
rect 339 220 342 222
rect 334 208 342 220
rect 344 208 349 224
rect 351 212 359 224
rect 351 210 354 212
rect 356 210 359 212
rect 351 208 359 210
rect 361 208 366 224
rect 368 222 375 224
rect 368 220 371 222
rect 373 220 375 222
rect 368 212 375 220
rect 401 217 406 224
rect 399 215 406 217
rect 399 213 401 215
rect 403 213 406 215
rect 368 208 374 212
rect 399 211 406 213
rect 334 206 339 208
rect 305 203 308 205
rect 310 203 312 205
rect 305 201 312 203
rect 305 196 310 201
rect 370 204 374 208
rect 401 206 406 211
rect 408 222 416 224
rect 408 220 411 222
rect 413 220 416 222
rect 408 208 416 220
rect 418 208 423 224
rect 425 212 433 224
rect 425 210 428 212
rect 430 210 433 212
rect 425 208 433 210
rect 435 208 440 224
rect 442 222 449 224
rect 442 220 445 222
rect 447 220 449 222
rect 442 212 449 220
rect 475 217 480 224
rect 473 215 480 217
rect 473 213 475 215
rect 477 213 480 215
rect 442 208 448 212
rect 473 211 480 213
rect 408 206 413 208
rect 370 196 376 204
rect 378 202 383 204
rect 378 200 385 202
rect 378 198 381 200
rect 383 198 385 200
rect 378 196 385 198
rect 444 204 448 208
rect 475 206 480 211
rect 482 222 490 224
rect 482 220 485 222
rect 487 220 490 222
rect 482 208 490 220
rect 492 208 497 224
rect 499 212 507 224
rect 499 210 502 212
rect 504 210 507 212
rect 499 208 507 210
rect 509 208 514 224
rect 516 222 523 224
rect 516 220 519 222
rect 521 220 523 222
rect 516 212 523 220
rect 516 208 522 212
rect 482 206 487 208
rect 444 196 450 204
rect 452 202 457 204
rect 452 200 459 202
rect 452 198 455 200
rect 457 198 459 200
rect 452 196 459 198
rect 518 204 522 208
rect 518 196 524 204
rect 526 202 531 204
rect 526 200 533 202
rect 526 198 529 200
rect 531 198 533 200
rect 526 196 533 198
rect -27 115 -22 120
rect -29 113 -22 115
rect -29 111 -27 113
rect -25 111 -22 113
rect -29 106 -22 111
rect -29 104 -27 106
rect -25 104 -22 106
rect -29 102 -22 104
rect -20 113 -12 120
rect 11 117 18 119
rect 11 115 13 117
rect 15 115 18 117
rect -20 102 -9 113
rect -18 96 -9 102
rect -18 94 -16 96
rect -14 94 -9 96
rect -18 92 -9 94
rect -7 92 -2 113
rect 0 105 5 113
rect 11 110 18 115
rect 11 108 13 110
rect 15 108 18 110
rect 11 106 18 108
rect 0 103 7 105
rect 0 101 3 103
rect 5 101 7 103
rect 13 101 18 106
rect 20 112 26 119
rect 59 117 66 119
rect 59 115 61 117
rect 63 115 66 117
rect 59 113 66 115
rect 20 105 28 112
rect 20 103 23 105
rect 25 103 28 105
rect 20 101 28 103
rect 0 99 7 101
rect 0 92 5 99
rect 22 99 28 101
rect 30 110 38 112
rect 30 108 33 110
rect 35 108 38 110
rect 30 103 38 108
rect 30 101 33 103
rect 35 101 38 103
rect 30 99 38 101
rect 40 103 47 112
rect 40 101 43 103
rect 45 101 47 103
rect 40 99 47 101
rect 61 92 66 113
rect 68 103 82 119
rect 68 101 71 103
rect 73 101 82 103
rect 84 117 92 119
rect 84 115 87 117
rect 89 115 92 117
rect 84 110 92 115
rect 84 108 87 110
rect 89 108 92 110
rect 84 101 92 108
rect 94 110 102 119
rect 94 108 97 110
rect 99 108 102 110
rect 94 101 102 108
rect 68 96 80 101
rect 68 94 71 96
rect 73 94 80 96
rect 68 92 80 94
rect 97 92 102 101
rect 104 104 109 119
rect 115 117 122 119
rect 115 115 117 117
rect 119 115 122 117
rect 115 110 122 115
rect 115 108 117 110
rect 119 108 122 110
rect 115 106 122 108
rect 104 102 111 104
rect 104 100 107 102
rect 109 100 111 102
rect 117 101 122 106
rect 124 112 130 119
rect 163 117 170 119
rect 163 115 165 117
rect 167 115 170 117
rect 163 113 170 115
rect 124 105 132 112
rect 124 103 127 105
rect 129 103 132 105
rect 124 101 132 103
rect 104 98 111 100
rect 104 92 109 98
rect 126 99 132 101
rect 134 110 142 112
rect 134 108 137 110
rect 139 108 142 110
rect 134 103 142 108
rect 134 101 137 103
rect 139 101 142 103
rect 134 99 142 101
rect 144 103 151 112
rect 144 101 147 103
rect 149 101 151 103
rect 144 99 151 101
rect 165 92 170 113
rect 172 103 186 119
rect 172 101 175 103
rect 177 101 186 103
rect 188 117 196 119
rect 188 115 191 117
rect 193 115 196 117
rect 188 110 196 115
rect 188 108 191 110
rect 193 108 196 110
rect 188 101 196 108
rect 198 110 206 119
rect 198 108 201 110
rect 203 108 206 110
rect 198 101 206 108
rect 172 96 184 101
rect 172 94 175 96
rect 177 94 184 96
rect 172 92 184 94
rect 201 92 206 101
rect 208 104 213 119
rect 249 112 255 119
rect 208 102 215 104
rect 208 100 211 102
rect 213 100 215 102
rect 208 98 215 100
rect 228 103 235 112
rect 228 101 230 103
rect 232 101 235 103
rect 228 99 235 101
rect 237 110 245 112
rect 237 108 240 110
rect 242 108 245 110
rect 237 103 245 108
rect 237 101 240 103
rect 242 101 245 103
rect 237 99 245 101
rect 247 105 255 112
rect 247 103 250 105
rect 252 103 255 105
rect 247 101 255 103
rect 257 117 264 119
rect 257 115 260 117
rect 262 115 264 117
rect 257 110 264 115
rect 295 113 303 120
rect 257 108 260 110
rect 262 108 264 110
rect 257 106 264 108
rect 257 101 262 106
rect 278 105 283 113
rect 276 103 283 105
rect 276 101 278 103
rect 280 101 283 103
rect 247 99 253 101
rect 208 92 213 98
rect 276 99 283 101
rect 278 92 283 99
rect 285 92 290 113
rect 292 102 303 113
rect 305 115 310 120
rect 305 113 312 115
rect 305 111 308 113
rect 310 111 312 113
rect 305 106 312 111
rect 305 104 308 106
rect 310 104 312 106
rect 327 105 332 110
rect 305 102 312 104
rect 325 103 332 105
rect 292 96 301 102
rect 325 101 327 103
rect 329 101 332 103
rect 325 99 332 101
rect 292 94 297 96
rect 299 94 301 96
rect 292 92 301 94
rect 327 92 332 99
rect 334 108 339 110
rect 370 112 376 120
rect 378 118 385 120
rect 378 116 381 118
rect 383 116 385 118
rect 378 114 385 116
rect 378 112 383 114
rect 370 108 374 112
rect 334 96 342 108
rect 334 94 337 96
rect 339 94 342 96
rect 334 92 342 94
rect 344 92 349 108
rect 351 106 359 108
rect 351 104 354 106
rect 356 104 359 106
rect 351 92 359 104
rect 361 92 366 108
rect 368 104 374 108
rect 401 105 406 110
rect 368 96 375 104
rect 399 103 406 105
rect 399 101 401 103
rect 403 101 406 103
rect 399 99 406 101
rect 368 94 371 96
rect 373 94 375 96
rect 368 92 375 94
rect 401 92 406 99
rect 408 108 413 110
rect 444 112 450 120
rect 452 118 459 120
rect 452 116 455 118
rect 457 116 459 118
rect 452 114 459 116
rect 452 112 457 114
rect 444 108 448 112
rect 408 96 416 108
rect 408 94 411 96
rect 413 94 416 96
rect 408 92 416 94
rect 418 92 423 108
rect 425 106 433 108
rect 425 104 428 106
rect 430 104 433 106
rect 425 92 433 104
rect 435 92 440 108
rect 442 104 448 108
rect 475 105 480 110
rect 442 96 449 104
rect 473 103 480 105
rect 473 101 475 103
rect 477 101 480 103
rect 473 99 480 101
rect 442 94 445 96
rect 447 94 449 96
rect 442 92 449 94
rect 475 92 480 99
rect 482 108 487 110
rect 518 112 524 120
rect 526 118 533 120
rect 526 116 529 118
rect 531 116 533 118
rect 526 114 533 116
rect 526 112 531 114
rect 518 108 522 112
rect 482 96 490 108
rect 482 94 485 96
rect 487 94 490 96
rect 482 92 490 94
rect 492 92 497 108
rect 499 106 507 108
rect 499 104 502 106
rect 504 104 507 106
rect 499 92 507 104
rect 509 92 514 108
rect 516 104 522 108
rect 516 96 523 104
rect 516 94 519 96
rect 521 94 523 96
rect 516 92 523 94
rect -18 78 -9 80
rect -18 76 -16 78
rect -14 76 -9 78
rect -29 70 -25 72
rect -18 70 -9 76
rect -29 68 -22 70
rect -29 66 -27 68
rect -25 66 -22 68
rect -29 61 -22 66
rect -29 59 -27 61
rect -25 59 -22 61
rect -29 57 -22 59
rect -27 52 -22 57
rect -20 59 -9 70
rect -7 59 -2 80
rect 0 73 5 80
rect 0 71 7 73
rect 22 71 28 73
rect 0 69 3 71
rect 5 69 7 71
rect 0 67 7 69
rect 0 59 5 67
rect 13 66 18 71
rect 11 64 18 66
rect 11 62 13 64
rect 15 62 18 64
rect -20 52 -12 59
rect 11 57 18 62
rect 11 55 13 57
rect 15 55 18 57
rect 11 53 18 55
rect 20 69 28 71
rect 20 67 23 69
rect 25 67 28 69
rect 20 60 28 67
rect 30 71 38 73
rect 30 69 33 71
rect 35 69 38 71
rect 30 64 38 69
rect 30 62 33 64
rect 35 62 38 64
rect 30 60 38 62
rect 40 71 47 73
rect 40 69 43 71
rect 45 69 47 71
rect 40 60 47 69
rect 20 53 26 60
rect 61 59 66 80
rect 59 57 66 59
rect 59 55 61 57
rect 63 55 66 57
rect 59 53 66 55
rect 68 78 80 80
rect 68 76 71 78
rect 73 76 80 78
rect 68 71 80 76
rect 97 71 102 80
rect 68 69 71 71
rect 73 69 82 71
rect 68 53 82 69
rect 84 64 92 71
rect 84 62 87 64
rect 89 62 92 64
rect 84 57 92 62
rect 84 55 87 57
rect 89 55 92 57
rect 84 53 92 55
rect 94 64 102 71
rect 94 62 97 64
rect 99 62 102 64
rect 94 53 102 62
rect 104 74 109 80
rect 104 72 111 74
rect 104 70 107 72
rect 109 70 111 72
rect 126 71 132 73
rect 104 68 111 70
rect 104 53 109 68
rect 117 66 122 71
rect 115 64 122 66
rect 115 62 117 64
rect 119 62 122 64
rect 115 57 122 62
rect 115 55 117 57
rect 119 55 122 57
rect 115 53 122 55
rect 124 69 132 71
rect 124 67 127 69
rect 129 67 132 69
rect 124 60 132 67
rect 134 71 142 73
rect 134 69 137 71
rect 139 69 142 71
rect 134 64 142 69
rect 134 62 137 64
rect 139 62 142 64
rect 134 60 142 62
rect 144 71 151 73
rect 144 69 147 71
rect 149 69 151 71
rect 144 60 151 69
rect 124 53 130 60
rect 165 59 170 80
rect 163 57 170 59
rect 163 55 165 57
rect 167 55 170 57
rect 163 53 170 55
rect 172 78 184 80
rect 172 76 175 78
rect 177 76 184 78
rect 172 71 184 76
rect 201 71 206 80
rect 172 69 175 71
rect 177 69 186 71
rect 172 53 186 69
rect 188 64 196 71
rect 188 62 191 64
rect 193 62 196 64
rect 188 57 196 62
rect 188 55 191 57
rect 193 55 196 57
rect 188 53 196 55
rect 198 64 206 71
rect 198 62 201 64
rect 203 62 206 64
rect 198 53 206 62
rect 208 74 213 80
rect 208 72 215 74
rect 208 70 211 72
rect 213 70 215 72
rect 208 68 215 70
rect 228 71 235 73
rect 228 69 230 71
rect 232 69 235 71
rect 208 53 213 68
rect 228 60 235 69
rect 237 71 245 73
rect 237 69 240 71
rect 242 69 245 71
rect 237 64 245 69
rect 237 62 240 64
rect 242 62 245 64
rect 237 60 245 62
rect 247 71 253 73
rect 278 73 283 80
rect 276 71 283 73
rect 247 69 255 71
rect 247 67 250 69
rect 252 67 255 69
rect 247 60 255 67
rect 249 53 255 60
rect 257 66 262 71
rect 276 69 278 71
rect 280 69 283 71
rect 276 67 283 69
rect 257 64 264 66
rect 257 62 260 64
rect 262 62 264 64
rect 257 57 264 62
rect 278 59 283 67
rect 285 59 290 80
rect 292 78 301 80
rect 292 76 297 78
rect 299 76 301 78
rect 292 70 301 76
rect 327 73 332 80
rect 325 71 332 73
rect 292 59 303 70
rect 257 55 260 57
rect 262 55 264 57
rect 257 53 264 55
rect 295 52 303 59
rect 305 68 312 70
rect 305 66 308 68
rect 310 66 312 68
rect 325 69 327 71
rect 329 69 332 71
rect 325 67 332 69
rect 305 61 312 66
rect 327 62 332 67
rect 334 78 342 80
rect 334 76 337 78
rect 339 76 342 78
rect 334 64 342 76
rect 344 64 349 80
rect 351 68 359 80
rect 351 66 354 68
rect 356 66 359 68
rect 351 64 359 66
rect 361 64 366 80
rect 368 78 375 80
rect 368 76 371 78
rect 373 76 375 78
rect 368 68 375 76
rect 401 73 406 80
rect 399 71 406 73
rect 399 69 401 71
rect 403 69 406 71
rect 368 64 374 68
rect 399 67 406 69
rect 334 62 339 64
rect 305 59 308 61
rect 310 59 312 61
rect 305 57 312 59
rect 305 52 310 57
rect 370 60 374 64
rect 401 62 406 67
rect 408 78 416 80
rect 408 76 411 78
rect 413 76 416 78
rect 408 64 416 76
rect 418 64 423 80
rect 425 68 433 80
rect 425 66 428 68
rect 430 66 433 68
rect 425 64 433 66
rect 435 64 440 80
rect 442 78 449 80
rect 442 76 445 78
rect 447 76 449 78
rect 442 68 449 76
rect 475 73 480 80
rect 473 71 480 73
rect 473 69 475 71
rect 477 69 480 71
rect 442 64 448 68
rect 473 67 480 69
rect 408 62 413 64
rect 370 52 376 60
rect 378 58 383 60
rect 378 56 385 58
rect 378 54 381 56
rect 383 54 385 56
rect 378 52 385 54
rect 444 60 448 64
rect 475 62 480 67
rect 482 78 490 80
rect 482 76 485 78
rect 487 76 490 78
rect 482 64 490 76
rect 492 64 497 80
rect 499 68 507 80
rect 499 66 502 68
rect 504 66 507 68
rect 499 64 507 66
rect 509 64 514 80
rect 516 78 523 80
rect 516 76 519 78
rect 521 76 523 78
rect 516 68 523 76
rect 516 64 522 68
rect 482 62 487 64
rect 444 52 450 60
rect 452 58 457 60
rect 452 56 459 58
rect 452 54 455 56
rect 457 54 459 56
rect 452 52 459 54
rect 518 60 522 64
rect 518 52 524 60
rect 526 58 531 60
rect 526 56 533 58
rect 526 54 529 56
rect 531 54 533 56
rect 526 52 533 54
<< alu1 >>
rect -33 297 537 302
rect -33 295 -26 297
rect -24 295 14 297
rect 16 295 24 297
rect 26 295 54 297
rect 56 295 107 297
rect 109 295 118 297
rect 120 295 128 297
rect 130 295 158 297
rect 160 295 211 297
rect 213 295 249 297
rect 251 295 259 297
rect 261 295 307 297
rect 309 295 537 297
rect -33 294 537 295
rect 11 285 23 289
rect 11 283 13 285
rect 15 283 23 285
rect 87 287 111 288
rect -29 280 -24 282
rect -29 278 -27 280
rect -25 278 -24 280
rect -29 276 -24 278
rect -29 257 -25 276
rect 3 272 7 281
rect -29 255 -27 257
rect -29 250 -25 255
rect -29 248 -27 250
rect -14 271 7 272
rect -14 269 -10 271
rect -8 269 4 271
rect 6 269 7 271
rect -14 268 7 269
rect -14 262 0 264
rect 2 262 7 264
rect -14 260 7 262
rect 3 258 7 260
rect 3 256 4 258
rect 6 256 7 258
rect 3 251 7 256
rect 11 263 15 283
rect 87 285 89 287
rect 91 285 111 287
rect 87 284 111 285
rect 35 280 40 281
rect 35 278 36 280
rect 38 278 40 280
rect 35 272 40 278
rect 11 261 16 263
rect 11 259 13 261
rect 15 259 16 261
rect 11 258 16 259
rect 11 256 12 258
rect 14 256 16 258
rect 11 254 16 256
rect 11 252 13 254
rect 15 252 16 254
rect 26 271 40 272
rect 26 269 30 271
rect 32 269 40 271
rect 26 268 40 269
rect 59 280 72 281
rect 59 278 61 280
rect 63 278 69 280
rect 71 278 72 280
rect 59 276 72 278
rect 59 275 69 276
rect 67 274 69 275
rect 71 274 72 276
rect 34 263 47 264
rect 34 261 40 263
rect 42 261 47 263
rect 34 260 47 261
rect 11 250 16 252
rect -29 244 -16 248
rect -29 243 -25 244
rect 43 256 47 260
rect 43 254 44 256
rect 46 254 47 256
rect 43 251 47 254
rect 51 263 56 265
rect 51 261 53 263
rect 55 261 56 263
rect 51 256 56 261
rect 67 267 72 274
rect 51 254 53 256
rect 55 254 56 256
rect 51 249 56 254
rect 51 243 63 249
rect 107 263 111 284
rect 107 261 108 263
rect 110 261 111 263
rect 107 256 111 261
rect 95 254 111 256
rect 95 252 97 254
rect 99 252 111 254
rect 95 251 111 252
rect 115 285 127 289
rect 115 283 117 285
rect 119 283 127 285
rect 191 287 215 288
rect 115 271 119 283
rect 191 285 193 287
rect 195 285 215 287
rect 191 284 215 285
rect 115 269 116 271
rect 118 269 119 271
rect 115 263 119 269
rect 139 280 144 281
rect 139 278 140 280
rect 142 278 144 280
rect 139 272 144 278
rect 115 261 120 263
rect 115 259 117 261
rect 119 259 120 261
rect 115 254 120 259
rect 115 252 117 254
rect 119 252 120 254
rect 130 271 144 272
rect 130 269 131 271
rect 133 269 134 271
rect 136 269 144 271
rect 130 268 144 269
rect 163 280 176 281
rect 163 278 165 280
rect 167 278 176 280
rect 163 276 176 278
rect 163 275 173 276
rect 171 274 173 275
rect 175 274 176 276
rect 138 263 151 264
rect 138 261 139 263
rect 141 261 144 263
rect 146 261 151 263
rect 138 260 151 261
rect 115 250 120 252
rect 147 256 151 260
rect 147 254 148 256
rect 150 254 151 256
rect 147 251 151 254
rect 155 263 160 265
rect 155 261 157 263
rect 159 261 160 263
rect 155 256 160 261
rect 171 267 176 274
rect 211 275 215 284
rect 211 273 212 275
rect 214 273 215 275
rect 155 254 157 256
rect 159 254 160 256
rect 155 249 160 254
rect 155 243 167 249
rect 211 256 215 273
rect 235 280 240 281
rect 235 278 237 280
rect 239 278 240 280
rect 235 272 240 278
rect 252 285 264 289
rect 252 283 260 285
rect 262 283 264 285
rect 235 271 249 272
rect 235 269 243 271
rect 245 269 249 271
rect 235 268 249 269
rect 199 254 215 256
rect 199 252 201 254
rect 203 252 215 254
rect 199 251 215 252
rect 228 263 241 264
rect 228 261 229 263
rect 231 261 233 263
rect 235 261 241 263
rect 228 260 241 261
rect 228 251 232 260
rect 260 266 264 283
rect 325 287 329 289
rect 325 285 330 287
rect 325 283 327 285
rect 329 283 330 285
rect 399 287 403 289
rect 276 280 280 281
rect 276 278 277 280
rect 279 278 280 280
rect 276 272 280 278
rect 276 271 297 272
rect 276 269 291 271
rect 293 269 297 271
rect 276 268 297 269
rect 307 280 312 282
rect 307 278 308 280
rect 310 278 312 280
rect 307 276 312 278
rect 260 264 261 266
rect 263 264 264 266
rect 260 263 264 264
rect 259 261 264 263
rect 259 259 260 261
rect 262 259 264 261
rect 259 254 264 259
rect 259 252 260 254
rect 262 252 264 254
rect 259 250 264 252
rect 276 263 281 264
rect 276 261 277 263
rect 279 262 281 263
rect 283 262 297 264
rect 279 261 297 262
rect 276 260 297 261
rect 276 251 280 260
rect 308 265 312 276
rect 308 263 309 265
rect 311 263 312 265
rect 308 257 312 263
rect 310 255 312 257
rect 308 250 312 255
rect 310 248 312 250
rect 299 244 312 248
rect 325 281 330 283
rect 325 273 329 281
rect 325 271 326 273
rect 328 271 329 273
rect 325 248 329 271
rect 334 265 336 267
rect 340 266 345 273
rect 340 264 341 266
rect 343 265 345 266
rect 343 264 353 265
rect 340 263 353 264
rect 340 261 341 263
rect 343 261 353 263
rect 340 259 353 261
rect 365 276 378 280
rect 365 274 368 276
rect 370 274 372 276
rect 365 273 372 274
rect 365 271 368 273
rect 370 271 372 273
rect 365 267 372 271
rect 370 260 372 262
rect 399 285 404 287
rect 399 283 401 285
rect 403 283 404 285
rect 473 287 477 289
rect 399 281 404 283
rect 399 269 403 281
rect 399 267 400 269
rect 402 267 403 269
rect 372 252 385 256
rect 380 251 385 252
rect 325 247 338 248
rect 380 249 381 251
rect 383 249 385 251
rect 325 245 327 247
rect 329 245 338 247
rect 325 244 338 245
rect 308 243 312 244
rect 380 243 385 249
rect 399 248 403 267
rect 415 271 421 273
rect 415 269 417 271
rect 419 269 421 271
rect 415 268 421 269
rect 408 265 410 267
rect 414 266 421 268
rect 414 264 415 266
rect 417 265 421 266
rect 417 264 427 265
rect 414 262 427 264
rect 415 259 427 262
rect 439 276 452 280
rect 439 271 445 276
rect 439 269 442 271
rect 444 269 445 271
rect 439 267 445 269
rect 444 260 446 262
rect 473 285 478 287
rect 473 283 475 285
rect 477 283 478 285
rect 473 281 478 283
rect 446 252 459 256
rect 454 251 459 252
rect 399 247 412 248
rect 454 249 455 251
rect 457 249 459 251
rect 399 245 401 247
rect 403 245 412 247
rect 399 244 412 245
rect 454 243 459 249
rect 473 248 477 281
rect 489 269 493 273
rect 482 265 484 267
rect 489 267 490 269
rect 492 267 493 269
rect 489 266 493 267
rect 491 265 493 266
rect 491 264 501 265
rect 489 259 501 264
rect 513 278 526 280
rect 513 276 516 278
rect 518 276 526 278
rect 513 271 519 276
rect 513 269 516 271
rect 518 269 519 271
rect 513 267 519 269
rect 518 260 520 262
rect 520 252 533 256
rect 528 251 533 252
rect 473 247 486 248
rect 528 249 529 251
rect 531 249 533 251
rect 473 245 475 247
rect 477 245 486 247
rect 473 244 486 245
rect 528 243 533 249
rect -33 237 537 238
rect -33 235 -26 237
rect -24 235 14 237
rect 16 235 87 237
rect 89 235 118 237
rect 120 235 191 237
rect 193 235 259 237
rect 261 235 307 237
rect 309 235 537 237
rect -33 225 537 235
rect -33 223 -26 225
rect -24 223 14 225
rect 16 223 87 225
rect 89 223 118 225
rect 120 223 191 225
rect 193 223 259 225
rect 261 223 307 225
rect 309 223 537 225
rect -33 222 537 223
rect -29 216 -25 217
rect -29 214 -28 216
rect -26 214 -16 216
rect -29 212 -16 214
rect -29 210 -27 212
rect -29 205 -25 210
rect -29 203 -27 205
rect -29 184 -25 203
rect 3 204 7 209
rect 3 202 4 204
rect 6 202 7 204
rect 3 200 7 202
rect -14 198 7 200
rect -14 196 0 198
rect 2 196 7 198
rect 11 208 16 210
rect 11 206 13 208
rect 15 206 16 208
rect 51 211 63 217
rect 11 204 16 206
rect 11 202 12 204
rect 14 202 16 204
rect 11 201 16 202
rect 11 199 13 201
rect 15 199 16 201
rect 11 197 16 199
rect 43 206 47 209
rect 43 204 44 206
rect 46 204 47 206
rect -29 182 -24 184
rect -29 180 -27 182
rect -25 180 -24 182
rect -29 178 -24 180
rect -14 191 7 192
rect -14 189 -10 191
rect -8 189 4 191
rect 6 189 7 191
rect -14 188 7 189
rect 3 179 7 188
rect 11 177 15 197
rect 43 200 47 204
rect 34 199 47 200
rect 34 197 40 199
rect 42 197 47 199
rect 34 196 47 197
rect 51 206 56 211
rect 51 204 53 206
rect 55 204 56 206
rect 51 199 56 204
rect 51 197 53 199
rect 55 197 56 199
rect 51 195 56 197
rect 26 191 40 192
rect 26 189 30 191
rect 32 189 40 191
rect 26 188 40 189
rect 11 175 13 177
rect 15 175 23 177
rect 11 171 23 175
rect 35 182 40 188
rect 35 180 36 182
rect 38 180 40 182
rect 35 179 40 180
rect 67 186 72 193
rect 95 208 111 209
rect 95 206 97 208
rect 99 206 111 208
rect 95 204 111 206
rect 107 199 111 204
rect 107 197 108 199
rect 110 197 111 199
rect 67 185 69 186
rect 59 184 69 185
rect 71 184 72 186
rect 59 182 72 184
rect 59 180 61 182
rect 63 180 72 182
rect 59 179 72 180
rect 107 176 111 197
rect 87 175 111 176
rect 87 173 89 175
rect 91 173 111 175
rect 87 172 111 173
rect 115 208 120 210
rect 115 206 117 208
rect 119 206 120 208
rect 155 211 167 217
rect 115 201 120 206
rect 115 199 117 201
rect 119 199 120 201
rect 115 197 120 199
rect 147 206 151 209
rect 147 204 148 206
rect 150 204 151 206
rect 115 191 119 197
rect 115 189 116 191
rect 118 189 119 191
rect 115 177 119 189
rect 147 200 151 204
rect 138 199 151 200
rect 138 197 139 199
rect 141 197 144 199
rect 146 197 151 199
rect 138 196 151 197
rect 155 206 160 211
rect 155 204 157 206
rect 159 204 160 206
rect 155 199 160 204
rect 155 197 157 199
rect 159 197 160 199
rect 155 195 160 197
rect 130 191 144 192
rect 130 189 131 191
rect 133 189 134 191
rect 136 189 144 191
rect 130 188 144 189
rect 115 175 117 177
rect 119 175 127 177
rect 115 171 127 175
rect 139 182 144 188
rect 139 180 140 182
rect 142 180 144 182
rect 139 179 144 180
rect 171 186 176 193
rect 199 208 215 209
rect 199 206 201 208
rect 203 206 215 208
rect 199 204 215 206
rect 171 185 173 186
rect 163 184 173 185
rect 175 184 176 186
rect 163 182 176 184
rect 163 180 165 182
rect 167 180 176 182
rect 163 179 176 180
rect 211 187 215 204
rect 228 200 232 209
rect 308 216 312 217
rect 299 212 312 216
rect 259 208 264 210
rect 228 199 241 200
rect 228 197 229 199
rect 231 197 233 199
rect 235 197 241 199
rect 228 196 241 197
rect 211 185 212 187
rect 214 185 215 187
rect 211 176 215 185
rect 235 191 249 192
rect 235 189 243 191
rect 245 189 249 191
rect 235 188 249 189
rect 259 206 260 208
rect 262 206 264 208
rect 259 201 264 206
rect 259 199 260 201
rect 262 199 264 201
rect 259 197 264 199
rect 235 182 240 188
rect 235 180 236 182
rect 238 180 240 182
rect 235 179 240 180
rect 260 196 264 197
rect 276 200 280 209
rect 276 199 297 200
rect 276 197 277 199
rect 279 198 297 199
rect 279 197 281 198
rect 276 196 281 197
rect 283 196 297 198
rect 260 194 261 196
rect 263 194 264 196
rect 260 177 264 194
rect 276 191 297 192
rect 276 189 291 191
rect 293 189 297 191
rect 276 188 297 189
rect 310 210 312 212
rect 308 205 312 210
rect 310 203 312 205
rect 276 182 280 188
rect 308 197 312 203
rect 308 195 309 197
rect 311 195 312 197
rect 308 184 312 195
rect 276 180 277 182
rect 279 180 280 182
rect 276 179 280 180
rect 307 182 312 184
rect 307 180 308 182
rect 310 180 312 182
rect 307 178 312 180
rect 325 215 338 216
rect 325 213 327 215
rect 329 213 338 215
rect 325 212 338 213
rect 325 189 329 212
rect 380 211 385 217
rect 380 209 381 211
rect 383 209 385 211
rect 325 187 326 189
rect 328 187 329 189
rect 380 208 385 209
rect 372 204 385 208
rect 399 215 412 216
rect 399 213 401 215
rect 403 213 412 215
rect 399 212 412 213
rect 334 193 336 195
rect 325 179 329 187
rect 340 199 353 201
rect 340 197 341 199
rect 343 197 353 199
rect 340 196 353 197
rect 340 194 341 196
rect 343 195 353 196
rect 370 198 372 200
rect 343 194 345 195
rect 340 187 345 194
rect 365 189 372 193
rect 365 187 368 189
rect 370 187 372 189
rect 365 186 372 187
rect 365 184 368 186
rect 370 184 372 186
rect 365 180 378 184
rect 191 175 215 176
rect 191 173 193 175
rect 195 173 215 175
rect 191 172 215 173
rect 252 175 260 177
rect 262 175 264 177
rect 252 171 264 175
rect 325 177 330 179
rect 325 175 327 177
rect 329 175 330 177
rect 325 173 330 175
rect 325 171 329 173
rect 399 193 403 212
rect 454 211 459 217
rect 454 209 455 211
rect 457 209 459 211
rect 399 191 400 193
rect 402 191 403 193
rect 399 179 403 191
rect 454 208 459 209
rect 446 204 459 208
rect 473 215 486 216
rect 473 213 475 215
rect 477 213 486 215
rect 473 212 486 213
rect 415 198 427 201
rect 408 193 410 195
rect 414 196 427 198
rect 414 194 415 196
rect 417 195 427 196
rect 444 198 446 200
rect 417 194 421 195
rect 414 192 421 194
rect 415 191 421 192
rect 415 189 417 191
rect 419 189 421 191
rect 415 187 421 189
rect 439 191 445 193
rect 439 189 442 191
rect 444 189 445 191
rect 439 184 445 189
rect 439 180 452 184
rect 399 177 404 179
rect 399 175 401 177
rect 403 175 404 177
rect 399 173 404 175
rect 399 171 403 173
rect 473 179 477 212
rect 528 211 533 217
rect 528 209 529 211
rect 531 209 533 211
rect 528 208 533 209
rect 520 204 533 208
rect 482 193 484 195
rect 489 196 501 201
rect 491 195 501 196
rect 518 198 520 200
rect 491 194 493 195
rect 489 193 493 194
rect 489 191 490 193
rect 492 191 493 193
rect 489 187 493 191
rect 513 191 519 193
rect 513 189 516 191
rect 518 189 519 191
rect 513 184 519 189
rect 513 182 516 184
rect 518 182 526 184
rect 513 180 526 182
rect 473 177 478 179
rect 473 175 475 177
rect 477 175 478 177
rect 473 173 478 175
rect 473 171 477 173
rect -33 165 537 166
rect -33 163 -26 165
rect -24 163 14 165
rect 16 163 24 165
rect 26 163 54 165
rect 56 163 107 165
rect 109 163 118 165
rect 120 163 128 165
rect 130 163 158 165
rect 160 163 211 165
rect 213 163 249 165
rect 251 163 259 165
rect 261 163 307 165
rect 309 163 537 165
rect -33 153 537 163
rect -33 151 -26 153
rect -24 151 14 153
rect 16 151 24 153
rect 26 151 54 153
rect 56 151 107 153
rect 109 151 118 153
rect 120 151 128 153
rect 130 151 158 153
rect 160 151 211 153
rect 213 151 249 153
rect 251 151 259 153
rect 261 151 307 153
rect 309 151 537 153
rect -33 150 537 151
rect 11 141 23 145
rect 11 139 13 141
rect 15 139 23 141
rect 87 143 111 144
rect -29 136 -24 138
rect -29 134 -27 136
rect -25 134 -24 136
rect -37 133 -24 134
rect -37 131 -36 133
rect -34 132 -24 133
rect -34 131 -25 132
rect -37 130 -25 131
rect -29 113 -25 130
rect 3 128 7 137
rect -29 111 -27 113
rect -29 106 -25 111
rect -29 104 -27 106
rect -14 127 7 128
rect -14 125 -10 127
rect -8 125 4 127
rect 6 125 7 127
rect -14 124 7 125
rect -14 118 0 120
rect 2 118 7 120
rect -14 116 7 118
rect 3 114 7 116
rect 3 112 4 114
rect 6 112 7 114
rect 3 107 7 112
rect 11 119 15 139
rect 87 141 89 143
rect 91 141 111 143
rect 87 140 111 141
rect 35 136 40 137
rect 35 134 36 136
rect 38 134 40 136
rect 35 128 40 134
rect 11 117 16 119
rect 11 115 13 117
rect 15 115 16 117
rect 11 114 16 115
rect 11 112 12 114
rect 14 112 16 114
rect 11 110 16 112
rect 11 108 13 110
rect 15 108 16 110
rect 26 127 40 128
rect 26 125 30 127
rect 32 125 40 127
rect 26 124 40 125
rect 59 136 72 137
rect 59 134 61 136
rect 63 134 69 136
rect 71 134 72 136
rect 59 132 72 134
rect 59 131 69 132
rect 67 130 69 131
rect 71 130 72 132
rect 34 119 47 120
rect 34 117 40 119
rect 42 117 44 119
rect 46 117 47 119
rect 34 116 47 117
rect 11 106 16 108
rect -29 100 -16 104
rect -29 99 -25 100
rect 43 111 47 116
rect 43 109 44 111
rect 46 109 47 111
rect 43 107 47 109
rect 51 119 56 121
rect 51 117 53 119
rect 55 117 56 119
rect 51 111 56 117
rect 67 123 72 130
rect 51 109 52 111
rect 54 109 56 111
rect 51 105 56 109
rect 51 99 63 105
rect 107 119 111 140
rect 107 117 108 119
rect 110 117 111 119
rect 107 112 111 117
rect 95 110 111 112
rect 95 108 97 110
rect 99 108 111 110
rect 95 107 111 108
rect 115 141 127 145
rect 115 139 117 141
rect 119 139 127 141
rect 191 143 215 144
rect 115 127 119 139
rect 191 141 193 143
rect 195 141 215 143
rect 191 140 215 141
rect 115 125 116 127
rect 118 125 119 127
rect 115 119 119 125
rect 139 136 144 137
rect 139 134 140 136
rect 142 134 144 136
rect 139 128 144 134
rect 115 117 120 119
rect 115 115 117 117
rect 119 115 120 117
rect 115 110 120 115
rect 115 108 117 110
rect 119 108 120 110
rect 130 127 144 128
rect 130 125 131 127
rect 133 125 134 127
rect 136 125 144 127
rect 130 124 144 125
rect 163 136 176 137
rect 163 134 165 136
rect 167 134 176 136
rect 163 132 176 134
rect 163 131 173 132
rect 171 130 173 131
rect 175 130 176 132
rect 138 119 151 120
rect 138 117 139 119
rect 141 117 144 119
rect 146 117 151 119
rect 138 116 151 117
rect 115 106 120 108
rect 147 112 151 116
rect 147 110 148 112
rect 150 110 151 112
rect 147 107 151 110
rect 155 119 160 121
rect 155 117 157 119
rect 159 117 160 119
rect 155 112 160 117
rect 171 123 176 130
rect 211 131 215 140
rect 211 129 212 131
rect 214 129 215 131
rect 155 110 157 112
rect 159 110 160 112
rect 155 105 160 110
rect 155 99 167 105
rect 211 112 215 129
rect 235 136 240 137
rect 235 134 237 136
rect 239 134 240 136
rect 235 128 240 134
rect 252 141 264 145
rect 252 139 260 141
rect 262 139 264 141
rect 235 127 249 128
rect 235 125 243 127
rect 245 125 249 127
rect 235 124 249 125
rect 199 110 215 112
rect 199 108 201 110
rect 203 108 215 110
rect 199 107 215 108
rect 228 119 241 120
rect 228 117 229 119
rect 231 117 233 119
rect 235 117 241 119
rect 228 116 241 117
rect 228 107 232 116
rect 260 122 264 139
rect 325 143 329 145
rect 325 141 330 143
rect 325 139 327 141
rect 329 139 330 141
rect 399 143 403 145
rect 276 136 280 137
rect 276 134 277 136
rect 279 134 280 136
rect 276 128 280 134
rect 276 127 297 128
rect 276 125 291 127
rect 293 125 297 127
rect 276 124 297 125
rect 307 136 312 138
rect 307 134 308 136
rect 310 134 312 136
rect 307 132 312 134
rect 260 120 261 122
rect 263 120 264 122
rect 260 119 264 120
rect 259 117 264 119
rect 259 115 260 117
rect 262 115 264 117
rect 259 110 264 115
rect 259 108 260 110
rect 262 108 264 110
rect 259 106 264 108
rect 276 119 281 120
rect 276 117 277 119
rect 279 118 281 119
rect 283 118 297 120
rect 279 117 297 118
rect 276 116 297 117
rect 276 107 280 116
rect 308 121 312 132
rect 308 119 309 121
rect 311 119 312 121
rect 308 113 312 119
rect 310 111 312 113
rect 308 106 312 111
rect 310 104 312 106
rect 299 100 312 104
rect 325 137 330 139
rect 325 129 329 137
rect 325 127 326 129
rect 328 127 329 129
rect 325 104 329 127
rect 334 121 336 123
rect 340 122 345 129
rect 340 120 341 122
rect 343 121 345 122
rect 343 120 353 121
rect 340 119 353 120
rect 340 117 341 119
rect 343 117 353 119
rect 340 115 353 117
rect 365 132 378 136
rect 365 130 368 132
rect 370 130 372 132
rect 365 129 372 130
rect 365 127 368 129
rect 370 127 372 129
rect 365 123 372 127
rect 370 116 372 118
rect 399 141 404 143
rect 399 139 401 141
rect 403 139 404 141
rect 473 143 477 145
rect 399 137 404 139
rect 399 125 403 137
rect 399 123 400 125
rect 402 123 403 125
rect 372 108 385 112
rect 380 107 385 108
rect 325 103 338 104
rect 380 105 381 107
rect 383 105 385 107
rect 325 101 327 103
rect 329 101 338 103
rect 325 100 338 101
rect 308 99 312 100
rect 380 99 385 105
rect 399 104 403 123
rect 415 127 421 129
rect 415 125 417 127
rect 419 125 421 127
rect 415 124 421 125
rect 408 121 410 123
rect 414 122 421 124
rect 414 120 415 122
rect 417 121 421 122
rect 417 120 427 121
rect 414 118 427 120
rect 415 115 427 118
rect 439 132 452 136
rect 439 127 445 132
rect 439 125 442 127
rect 444 125 445 127
rect 439 123 445 125
rect 444 116 446 118
rect 473 141 478 143
rect 473 139 475 141
rect 477 139 478 141
rect 473 137 478 139
rect 446 108 459 112
rect 454 107 459 108
rect 399 103 412 104
rect 454 105 455 107
rect 457 105 459 107
rect 399 101 401 103
rect 403 101 412 103
rect 399 100 412 101
rect 454 99 459 105
rect 473 104 477 137
rect 489 125 493 129
rect 482 121 484 123
rect 489 123 490 125
rect 492 123 493 125
rect 489 122 493 123
rect 491 121 493 122
rect 491 120 501 121
rect 489 115 501 120
rect 513 134 526 136
rect 513 132 516 134
rect 518 132 526 134
rect 513 127 519 132
rect 513 125 516 127
rect 518 125 519 127
rect 513 123 519 125
rect 518 116 520 118
rect 520 108 533 112
rect 528 107 533 108
rect 473 103 486 104
rect 528 105 529 107
rect 531 105 533 107
rect 473 101 475 103
rect 477 101 486 103
rect 473 100 486 101
rect 528 99 533 105
rect -33 93 537 94
rect -33 91 -26 93
rect -24 91 14 93
rect 16 91 87 93
rect 89 91 118 93
rect 120 91 191 93
rect 193 91 259 93
rect 261 91 307 93
rect 309 91 537 93
rect -33 81 537 91
rect -33 79 -26 81
rect -24 79 14 81
rect 16 79 87 81
rect 89 79 118 81
rect 120 79 191 81
rect 193 79 259 81
rect 261 79 307 81
rect 309 79 537 81
rect -33 78 537 79
rect -29 68 -16 72
rect -29 66 -27 68
rect -29 61 -25 66
rect -29 59 -27 61
rect -29 49 -25 59
rect 3 60 7 65
rect -29 47 -28 49
rect -26 47 -25 49
rect -29 40 -25 47
rect 3 58 4 60
rect 6 58 7 60
rect 3 56 7 58
rect -14 54 7 56
rect -14 52 0 54
rect 2 52 7 54
rect 11 64 16 66
rect 11 62 13 64
rect 15 62 16 64
rect 51 67 63 73
rect 11 60 16 62
rect 11 58 12 60
rect 14 58 16 60
rect 11 57 16 58
rect 11 55 13 57
rect 15 55 16 57
rect 11 53 16 55
rect 43 62 47 65
rect 43 60 44 62
rect 46 60 47 62
rect -29 38 -24 40
rect -29 36 -27 38
rect -25 36 -24 38
rect -29 34 -24 36
rect -14 47 7 48
rect -14 45 -10 47
rect -8 45 4 47
rect 6 45 7 47
rect -14 44 7 45
rect 3 35 7 44
rect 11 33 15 53
rect 43 56 47 60
rect 34 55 47 56
rect 34 53 40 55
rect 42 53 47 55
rect 34 52 47 53
rect 51 62 56 67
rect 51 60 53 62
rect 55 60 56 62
rect 51 55 56 60
rect 51 53 53 55
rect 55 53 56 55
rect 51 51 56 53
rect 26 47 40 48
rect 26 45 30 47
rect 32 45 40 47
rect 26 44 40 45
rect 11 31 13 33
rect 15 31 23 33
rect 11 27 23 31
rect 35 38 40 44
rect 35 36 36 38
rect 38 36 40 38
rect 35 35 40 36
rect 67 42 72 49
rect 95 64 111 65
rect 95 62 97 64
rect 99 62 111 64
rect 95 60 111 62
rect 107 55 111 60
rect 107 53 108 55
rect 110 53 111 55
rect 67 41 69 42
rect 59 40 69 41
rect 71 40 72 42
rect 59 38 72 40
rect 59 36 61 38
rect 63 36 72 38
rect 59 35 72 36
rect 107 32 111 53
rect 87 31 111 32
rect 87 29 89 31
rect 91 29 111 31
rect 87 28 111 29
rect 115 64 120 66
rect 115 62 117 64
rect 119 62 120 64
rect 155 67 167 73
rect 115 57 120 62
rect 115 55 117 57
rect 119 55 120 57
rect 115 53 120 55
rect 147 62 151 65
rect 147 60 148 62
rect 150 60 151 62
rect 115 47 119 53
rect 115 45 116 47
rect 118 45 119 47
rect 115 33 119 45
rect 147 56 151 60
rect 138 55 151 56
rect 138 53 139 55
rect 141 53 144 55
rect 146 53 151 55
rect 138 52 151 53
rect 155 62 160 67
rect 155 60 157 62
rect 159 60 160 62
rect 155 55 160 60
rect 155 53 157 55
rect 159 53 160 55
rect 155 51 160 53
rect 130 47 144 48
rect 130 45 134 47
rect 136 45 144 47
rect 130 44 144 45
rect 115 31 117 33
rect 119 31 127 33
rect 115 27 127 31
rect 139 38 144 44
rect 139 36 140 38
rect 142 36 144 38
rect 139 35 144 36
rect 171 42 176 49
rect 199 64 215 65
rect 199 62 201 64
rect 203 62 215 64
rect 199 60 215 62
rect 171 41 173 42
rect 163 40 173 41
rect 175 40 176 42
rect 163 38 176 40
rect 163 36 165 38
rect 167 36 176 38
rect 163 35 176 36
rect 211 43 215 60
rect 228 63 232 65
rect 228 61 229 63
rect 231 61 232 63
rect 228 56 232 61
rect 308 72 312 73
rect 299 68 312 72
rect 259 64 264 66
rect 228 55 241 56
rect 228 53 233 55
rect 235 53 241 55
rect 228 52 241 53
rect 211 41 212 43
rect 214 41 215 43
rect 211 32 215 41
rect 235 47 249 48
rect 235 45 237 47
rect 239 45 243 47
rect 245 45 249 47
rect 235 44 249 45
rect 259 62 260 64
rect 262 62 264 64
rect 259 57 264 62
rect 259 55 260 57
rect 262 55 264 57
rect 259 53 264 55
rect 235 35 240 44
rect 260 52 264 53
rect 276 63 280 65
rect 276 61 277 63
rect 279 61 280 63
rect 276 56 280 61
rect 276 54 297 56
rect 276 52 281 54
rect 283 52 297 54
rect 260 50 261 52
rect 263 50 264 52
rect 260 33 264 50
rect 276 47 297 48
rect 276 45 277 47
rect 279 45 291 47
rect 293 45 297 47
rect 276 44 297 45
rect 310 66 312 68
rect 308 61 312 66
rect 310 59 312 61
rect 276 35 280 44
rect 308 53 312 59
rect 308 51 309 53
rect 311 51 312 53
rect 308 40 312 51
rect 307 38 312 40
rect 307 36 308 38
rect 310 36 312 38
rect 307 34 312 36
rect 325 71 338 72
rect 325 69 327 71
rect 329 69 338 71
rect 325 68 338 69
rect 325 45 329 68
rect 380 67 385 73
rect 380 65 381 67
rect 383 65 385 67
rect 325 43 326 45
rect 328 43 329 45
rect 380 64 385 65
rect 372 60 385 64
rect 399 71 412 72
rect 399 69 401 71
rect 403 69 412 71
rect 399 68 412 69
rect 334 49 336 51
rect 325 35 329 43
rect 340 55 353 57
rect 340 53 341 55
rect 343 53 353 55
rect 340 52 353 53
rect 340 50 341 52
rect 343 51 353 52
rect 370 54 372 56
rect 343 50 345 51
rect 340 43 345 50
rect 365 45 372 49
rect 365 43 368 45
rect 370 43 372 45
rect 365 42 372 43
rect 365 40 368 42
rect 370 40 372 42
rect 365 36 378 40
rect 191 31 215 32
rect 191 29 193 31
rect 195 29 215 31
rect 191 28 215 29
rect 252 31 260 33
rect 262 31 264 33
rect 252 27 264 31
rect 325 33 330 35
rect 325 31 327 33
rect 329 31 330 33
rect 325 29 330 31
rect 325 27 329 29
rect 399 49 403 68
rect 454 67 459 73
rect 454 65 455 67
rect 457 65 459 67
rect 399 47 400 49
rect 402 47 403 49
rect 399 35 403 47
rect 454 64 459 65
rect 446 60 459 64
rect 473 71 486 72
rect 473 69 475 71
rect 477 69 486 71
rect 473 68 486 69
rect 415 54 427 57
rect 408 49 410 51
rect 414 52 427 54
rect 414 50 415 52
rect 417 51 427 52
rect 444 54 446 56
rect 417 50 421 51
rect 414 48 421 50
rect 415 47 421 48
rect 415 45 417 47
rect 419 45 421 47
rect 415 43 421 45
rect 439 47 445 49
rect 439 45 442 47
rect 444 45 445 47
rect 439 40 445 45
rect 439 36 452 40
rect 399 33 404 35
rect 399 31 401 33
rect 403 31 404 33
rect 399 29 404 31
rect 399 27 403 29
rect 473 35 477 68
rect 528 67 533 73
rect 528 65 529 67
rect 531 65 533 67
rect 528 64 533 65
rect 520 60 533 64
rect 482 49 484 51
rect 489 52 501 57
rect 491 51 501 52
rect 518 54 520 56
rect 491 50 493 51
rect 489 49 493 50
rect 489 47 490 49
rect 492 47 493 49
rect 489 43 493 47
rect 513 47 519 49
rect 513 45 516 47
rect 518 45 519 47
rect 513 40 519 45
rect 513 38 516 40
rect 518 38 526 40
rect 513 36 526 38
rect 473 33 478 35
rect 473 31 475 33
rect 477 31 478 33
rect 473 29 478 31
rect 473 27 477 29
rect -33 21 537 22
rect -33 19 -26 21
rect -24 19 14 21
rect 16 19 24 21
rect 26 19 54 21
rect 56 19 107 21
rect 109 19 118 21
rect 120 19 128 21
rect 130 19 158 21
rect 160 19 211 21
rect 213 19 249 21
rect 251 19 259 21
rect 261 19 307 21
rect 309 19 537 21
rect -33 14 537 19
<< alu2 >>
rect 321 296 493 300
rect 35 280 72 281
rect 35 278 36 280
rect 38 278 61 280
rect 63 278 69 280
rect 71 278 72 280
rect 35 277 72 278
rect 139 280 171 281
rect 139 278 140 280
rect 142 278 165 280
rect 167 278 171 280
rect 35 276 67 277
rect 139 276 171 278
rect 236 280 240 281
rect 236 278 237 280
rect 239 278 240 280
rect 236 277 240 278
rect 276 280 280 281
rect 276 278 277 280
rect 279 278 280 280
rect 276 277 280 278
rect 211 275 224 276
rect 211 273 212 275
rect 214 273 224 275
rect 211 272 224 273
rect 3 271 119 272
rect 3 269 4 271
rect 6 269 116 271
rect 118 269 119 271
rect 3 268 119 269
rect 130 271 134 272
rect 130 269 131 271
rect 133 269 134 271
rect 130 268 134 269
rect 107 263 142 264
rect 107 261 108 263
rect 110 261 139 263
rect 141 261 142 263
rect 107 260 142 261
rect 3 258 16 259
rect 3 256 4 258
rect 6 256 12 258
rect 14 256 16 258
rect 3 254 16 256
rect 43 256 56 257
rect 43 254 44 256
rect 46 254 53 256
rect 55 254 56 256
rect 43 253 56 254
rect 147 256 160 257
rect 147 254 148 256
rect 150 254 157 256
rect 159 254 160 256
rect 147 253 160 254
rect 220 243 224 272
rect 321 274 325 296
rect 383 285 420 289
rect 321 273 329 274
rect 321 271 326 273
rect 328 271 329 273
rect 321 270 329 271
rect 367 273 371 276
rect 367 271 368 273
rect 370 271 371 273
rect 260 266 269 267
rect 340 266 344 267
rect 260 264 261 266
rect 263 264 269 266
rect 308 265 345 266
rect 228 263 232 264
rect 260 263 269 264
rect 228 261 229 263
rect 231 261 232 263
rect 228 260 232 261
rect 264 255 269 263
rect 276 263 280 264
rect 276 261 277 263
rect 279 261 280 263
rect 308 263 309 265
rect 311 263 345 265
rect 308 262 341 263
rect 276 260 280 261
rect 340 261 341 262
rect 343 261 345 263
rect 340 259 345 261
rect 367 255 371 271
rect 264 251 371 255
rect 383 243 387 285
rect 416 271 420 285
rect 220 239 387 243
rect 393 269 403 270
rect 393 267 400 269
rect 402 267 403 269
rect 393 266 403 267
rect 416 269 417 271
rect 419 269 420 271
rect 393 236 397 266
rect 416 263 420 269
rect 489 269 493 296
rect 489 267 490 269
rect 492 267 493 269
rect 489 262 493 267
rect 515 278 519 279
rect 515 276 516 278
rect 518 276 519 278
rect 515 236 519 276
rect 393 232 519 236
rect 393 224 519 228
rect 220 217 387 221
rect -29 216 -25 217
rect -29 214 -28 216
rect -26 214 -25 216
rect -29 213 -25 214
rect 43 206 56 207
rect 3 204 16 206
rect 3 202 4 204
rect 6 202 12 204
rect 14 202 16 204
rect 43 204 44 206
rect 46 204 53 206
rect 55 204 56 206
rect 43 203 56 204
rect 147 206 160 207
rect 147 204 148 206
rect 150 204 157 206
rect 159 204 160 206
rect 147 203 160 204
rect 3 201 16 202
rect 107 199 142 200
rect 107 197 108 199
rect 110 197 139 199
rect 141 197 142 199
rect 107 196 142 197
rect 3 191 119 192
rect 3 189 4 191
rect 6 189 116 191
rect 118 189 119 191
rect 3 188 119 189
rect 130 191 134 192
rect 130 189 131 191
rect 133 189 134 191
rect 130 188 134 189
rect 220 188 224 217
rect 264 205 371 209
rect 228 199 232 200
rect 228 197 229 199
rect 231 197 232 199
rect 264 197 269 205
rect 228 196 232 197
rect 260 196 269 197
rect 276 199 280 200
rect 276 197 277 199
rect 279 197 280 199
rect 340 199 345 201
rect 340 198 341 199
rect 276 196 280 197
rect 308 197 341 198
rect 343 197 345 199
rect 260 194 261 196
rect 263 194 269 196
rect 308 195 309 197
rect 311 195 345 197
rect 308 194 345 195
rect 260 193 269 194
rect 340 193 344 194
rect 211 187 224 188
rect 211 185 212 187
rect 214 185 224 187
rect 211 184 224 185
rect 321 189 329 190
rect 321 187 326 189
rect 328 187 329 189
rect 321 186 329 187
rect 367 189 371 205
rect 367 187 368 189
rect 370 187 371 189
rect 35 182 67 184
rect 35 180 36 182
rect 38 180 61 182
rect 63 180 67 182
rect 35 179 67 180
rect 139 182 171 184
rect 139 180 140 182
rect 142 180 165 182
rect 167 180 171 182
rect 139 179 171 180
rect 235 182 239 183
rect 235 180 236 182
rect 238 180 239 182
rect 235 179 239 180
rect 276 182 280 183
rect 276 180 277 182
rect 279 180 280 182
rect 276 179 280 180
rect 321 164 325 186
rect 367 184 371 187
rect 383 175 387 217
rect 393 194 397 224
rect 393 193 403 194
rect 393 191 400 193
rect 402 191 403 193
rect 393 190 403 191
rect 416 191 420 197
rect 416 189 417 191
rect 419 189 420 191
rect 416 175 420 189
rect 383 171 420 175
rect 489 193 493 198
rect 489 191 490 193
rect 492 191 493 193
rect 489 164 493 191
rect 515 184 519 224
rect 515 182 516 184
rect 518 182 519 184
rect 515 181 519 182
rect 321 160 493 164
rect 321 152 493 156
rect -37 147 -33 148
rect -37 145 -36 147
rect -34 145 -33 147
rect -37 133 -33 145
rect -37 131 -36 133
rect -34 131 -33 133
rect 35 136 72 137
rect 35 134 36 136
rect 38 134 61 136
rect 63 134 69 136
rect 71 134 72 136
rect 35 132 72 134
rect 139 136 171 137
rect 139 134 140 136
rect 142 134 165 136
rect 167 134 171 136
rect 139 132 171 134
rect 235 136 240 137
rect 235 134 237 136
rect 239 134 240 136
rect 235 133 240 134
rect 276 136 280 137
rect 276 134 277 136
rect 279 134 280 136
rect 276 133 280 134
rect -37 130 -33 131
rect 211 131 224 132
rect 211 129 212 131
rect 214 129 224 131
rect 211 128 224 129
rect 3 127 119 128
rect 3 125 4 127
rect 6 125 116 127
rect 118 125 119 127
rect 3 124 119 125
rect 130 127 134 128
rect 130 125 131 127
rect 133 125 134 127
rect 130 124 134 125
rect 43 119 56 120
rect 43 117 44 119
rect 46 117 56 119
rect 43 116 56 117
rect 107 119 142 120
rect 107 117 108 119
rect 110 117 139 119
rect 141 117 142 119
rect 107 116 142 117
rect 3 114 16 115
rect 3 112 4 114
rect 6 112 12 114
rect 14 112 16 114
rect 147 112 160 113
rect 3 110 16 112
rect 43 111 56 112
rect 43 109 44 111
rect 46 109 52 111
rect 54 109 56 111
rect 147 110 148 112
rect 150 110 157 112
rect 159 110 160 112
rect 147 109 160 110
rect 43 108 56 109
rect 220 99 224 128
rect 321 130 325 152
rect 383 141 420 145
rect 321 129 329 130
rect 321 127 326 129
rect 328 127 329 129
rect 321 126 329 127
rect 367 129 371 132
rect 367 127 368 129
rect 370 127 371 129
rect 260 122 269 123
rect 340 122 344 123
rect 260 120 261 122
rect 263 120 269 122
rect 308 121 345 122
rect 228 119 232 120
rect 260 119 269 120
rect 228 117 229 119
rect 231 117 232 119
rect 228 116 232 117
rect 264 111 269 119
rect 276 119 280 120
rect 276 117 277 119
rect 279 117 280 119
rect 308 119 309 121
rect 311 119 345 121
rect 308 118 341 119
rect 276 116 280 117
rect 340 117 341 118
rect 343 117 345 119
rect 340 115 345 117
rect 367 111 371 127
rect 264 107 371 111
rect 383 99 387 141
rect 416 127 420 141
rect 220 95 387 99
rect 393 125 403 126
rect 393 123 400 125
rect 402 123 403 125
rect 393 122 403 123
rect 416 125 417 127
rect 419 125 420 127
rect 393 92 397 122
rect 416 119 420 125
rect 489 125 493 152
rect 489 123 490 125
rect 492 123 493 125
rect 489 118 493 123
rect 515 134 519 135
rect 515 132 516 134
rect 518 132 519 134
rect 515 92 519 132
rect 393 88 519 92
rect 393 80 519 84
rect 220 73 387 77
rect 43 62 56 63
rect 3 60 16 62
rect 3 58 4 60
rect 6 58 12 60
rect 14 58 16 60
rect 43 60 44 62
rect 46 60 53 62
rect 55 60 56 62
rect 43 59 56 60
rect 147 62 160 63
rect 147 60 148 62
rect 150 60 157 62
rect 159 60 160 62
rect 147 59 160 60
rect 3 57 16 58
rect 107 55 142 56
rect 107 53 108 55
rect 110 53 139 55
rect 141 53 142 55
rect 107 52 142 53
rect -29 49 -25 50
rect -29 47 -28 49
rect -26 47 -25 49
rect -29 46 -25 47
rect 3 47 119 48
rect 3 45 4 47
rect 6 45 116 47
rect 118 45 119 47
rect 3 44 119 45
rect 220 44 224 73
rect 228 63 232 64
rect 228 61 229 63
rect 231 61 232 63
rect 228 59 232 61
rect 264 63 371 65
rect 264 61 277 63
rect 279 61 371 63
rect 264 53 269 61
rect 276 60 280 61
rect 340 55 345 57
rect 340 54 341 55
rect 260 52 269 53
rect 260 50 261 52
rect 263 50 269 52
rect 308 53 341 54
rect 343 53 345 55
rect 308 51 309 53
rect 311 51 345 53
rect 308 50 345 51
rect 260 49 269 50
rect 340 49 344 50
rect 236 47 240 48
rect 236 45 237 47
rect 239 45 240 47
rect 236 44 240 45
rect 276 47 280 48
rect 276 45 277 47
rect 279 45 280 47
rect 276 44 280 45
rect 321 45 329 46
rect 211 43 224 44
rect 211 41 212 43
rect 214 41 224 43
rect 211 40 224 41
rect 321 43 326 45
rect 328 43 329 45
rect 321 42 329 43
rect 367 45 371 61
rect 367 43 368 45
rect 370 43 371 45
rect 35 38 67 40
rect 35 36 36 38
rect 38 36 61 38
rect 63 36 67 38
rect 35 35 67 36
rect 139 38 171 40
rect 139 36 140 38
rect 142 36 165 38
rect 167 36 171 38
rect 139 35 171 36
rect 321 20 325 42
rect 367 40 371 43
rect 383 31 387 73
rect 393 50 397 80
rect 393 49 403 50
rect 393 47 400 49
rect 402 47 403 49
rect 393 46 403 47
rect 416 47 420 53
rect 416 45 417 47
rect 419 45 420 47
rect 416 31 420 45
rect 383 27 420 31
rect 489 49 493 54
rect 489 47 490 49
rect 492 47 493 49
rect 489 20 493 47
rect 515 40 519 80
rect 515 38 516 40
rect 518 38 519 40
rect 515 37 519 38
rect 321 16 493 20
<< alu3 >>
rect 67 280 280 281
rect 67 278 69 280
rect 71 278 237 280
rect 239 278 277 280
rect 279 278 280 280
rect 67 277 280 278
rect -29 271 136 272
rect -29 269 131 271
rect 133 269 136 271
rect -29 268 136 269
rect -29 216 -25 268
rect 51 263 280 264
rect 51 261 229 263
rect 231 261 277 263
rect 279 261 280 263
rect 51 260 280 261
rect 51 256 56 260
rect 51 254 53 256
rect 55 254 56 256
rect 51 253 56 254
rect -29 214 -28 216
rect -26 214 -25 216
rect -29 210 -25 214
rect 51 206 232 207
rect 51 204 53 206
rect 55 204 232 206
rect 51 203 232 204
rect 228 200 232 203
rect 228 199 280 200
rect 228 197 229 199
rect 231 197 277 199
rect 279 197 280 199
rect 228 196 280 197
rect 132 192 136 193
rect -29 191 136 192
rect -29 189 131 191
rect 133 189 136 191
rect -29 188 136 189
rect -29 148 -25 188
rect 60 182 280 183
rect 60 180 61 182
rect 63 180 236 182
rect 238 180 277 182
rect 279 180 280 182
rect 60 179 280 180
rect -37 147 -25 148
rect -37 145 -36 147
rect -34 145 -25 147
rect -37 144 -25 145
rect -29 132 -25 144
rect 68 136 280 137
rect 68 134 69 136
rect 71 134 237 136
rect 239 134 277 136
rect 279 134 280 136
rect 68 133 280 134
rect -29 127 136 128
rect -29 125 131 127
rect 133 125 136 127
rect -29 124 136 125
rect -29 49 -25 124
rect 42 119 280 120
rect 42 117 44 119
rect 46 117 229 119
rect 231 117 277 119
rect 279 117 280 119
rect 42 116 280 117
rect 43 63 280 64
rect 43 62 229 63
rect 43 60 44 62
rect 46 61 229 62
rect 231 61 277 63
rect 279 61 280 63
rect 46 60 280 61
rect 43 59 280 60
rect -29 47 -28 49
rect -26 47 -25 49
rect -29 46 -25 47
rect 78 44 88 48
rect 235 47 280 48
rect 235 45 237 47
rect 239 45 277 47
rect 279 45 280 47
rect 235 44 280 45
<< ptie >>
rect -28 297 -22 299
rect -28 295 -26 297
rect -24 295 -22 297
rect 12 297 18 299
rect 12 295 14 297
rect 16 295 18 297
rect -28 293 -22 295
rect 12 293 18 295
rect 52 297 58 299
rect 52 295 54 297
rect 56 295 58 297
rect 52 293 58 295
rect 116 297 122 299
rect 116 295 118 297
rect 120 295 122 297
rect 116 293 122 295
rect 156 297 162 299
rect 156 295 158 297
rect 160 295 162 297
rect 156 293 162 295
rect 257 297 263 299
rect 257 295 259 297
rect 261 295 263 297
rect 305 297 311 299
rect 305 295 307 297
rect 309 295 311 297
rect 257 293 263 295
rect 305 293 311 295
rect -28 165 -22 167
rect 12 165 18 167
rect -28 163 -26 165
rect -24 163 -22 165
rect -28 161 -22 163
rect 12 163 14 165
rect 16 163 18 165
rect 12 161 18 163
rect 52 165 58 167
rect 52 163 54 165
rect 56 163 58 165
rect 52 161 58 163
rect 116 165 122 167
rect 116 163 118 165
rect 120 163 122 165
rect 116 161 122 163
rect 156 165 162 167
rect 156 163 158 165
rect 160 163 162 165
rect 156 161 162 163
rect 257 165 263 167
rect 305 165 311 167
rect 257 163 259 165
rect 261 163 263 165
rect 257 161 263 163
rect 305 163 307 165
rect 309 163 311 165
rect 305 161 311 163
rect -28 153 -22 155
rect -28 151 -26 153
rect -24 151 -22 153
rect 12 153 18 155
rect 12 151 14 153
rect 16 151 18 153
rect -28 149 -22 151
rect 12 149 18 151
rect 52 153 58 155
rect 52 151 54 153
rect 56 151 58 153
rect 52 149 58 151
rect 116 153 122 155
rect 116 151 118 153
rect 120 151 122 153
rect 116 149 122 151
rect 156 153 162 155
rect 156 151 158 153
rect 160 151 162 153
rect 156 149 162 151
rect 257 153 263 155
rect 257 151 259 153
rect 261 151 263 153
rect 305 153 311 155
rect 305 151 307 153
rect 309 151 311 153
rect 257 149 263 151
rect 305 149 311 151
rect -28 21 -22 23
rect 12 21 18 23
rect -28 19 -26 21
rect -24 19 -22 21
rect -28 17 -22 19
rect 12 19 14 21
rect 16 19 18 21
rect 12 17 18 19
rect 52 21 58 23
rect 52 19 54 21
rect 56 19 58 21
rect 52 17 58 19
rect 116 21 122 23
rect 116 19 118 21
rect 120 19 122 21
rect 116 17 122 19
rect 156 21 162 23
rect 156 19 158 21
rect 160 19 162 21
rect 156 17 162 19
rect 257 21 263 23
rect 305 21 311 23
rect 257 19 259 21
rect 261 19 263 21
rect 257 17 263 19
rect 305 19 307 21
rect 309 19 311 21
rect 305 17 311 19
<< ntie >>
rect -28 237 -22 239
rect -28 235 -26 237
rect -24 235 -22 237
rect 12 237 18 239
rect -28 233 -22 235
rect 12 235 14 237
rect 16 235 18 237
rect 85 237 91 239
rect 12 233 18 235
rect 85 235 87 237
rect 89 235 91 237
rect 116 237 122 239
rect 85 233 91 235
rect 116 235 118 237
rect 120 235 122 237
rect 189 237 195 239
rect 116 233 122 235
rect 189 235 191 237
rect 193 235 195 237
rect 257 237 263 239
rect 189 233 195 235
rect 257 235 259 237
rect 261 235 263 237
rect 305 237 311 239
rect 257 233 263 235
rect 305 235 307 237
rect 309 235 311 237
rect 305 233 311 235
rect -28 225 -22 227
rect -28 223 -26 225
rect -24 223 -22 225
rect 12 225 18 227
rect -28 221 -22 223
rect 12 223 14 225
rect 16 223 18 225
rect 85 225 91 227
rect 12 221 18 223
rect 85 223 87 225
rect 89 223 91 225
rect 116 225 122 227
rect 85 221 91 223
rect 116 223 118 225
rect 120 223 122 225
rect 189 225 195 227
rect 116 221 122 223
rect 189 223 191 225
rect 193 223 195 225
rect 257 225 263 227
rect 189 221 195 223
rect 257 223 259 225
rect 261 223 263 225
rect 305 225 311 227
rect 257 221 263 223
rect 305 223 307 225
rect 309 223 311 225
rect 305 221 311 223
rect -28 93 -22 95
rect -28 91 -26 93
rect -24 91 -22 93
rect 12 93 18 95
rect -28 89 -22 91
rect 12 91 14 93
rect 16 91 18 93
rect 85 93 91 95
rect 12 89 18 91
rect 85 91 87 93
rect 89 91 91 93
rect 116 93 122 95
rect 85 89 91 91
rect 116 91 118 93
rect 120 91 122 93
rect 189 93 195 95
rect 116 89 122 91
rect 189 91 191 93
rect 193 91 195 93
rect 257 93 263 95
rect 189 89 195 91
rect 257 91 259 93
rect 261 91 263 93
rect 305 93 311 95
rect 257 89 263 91
rect 305 91 307 93
rect 309 91 311 93
rect 305 89 311 91
rect -28 81 -22 83
rect -28 79 -26 81
rect -24 79 -22 81
rect 12 81 18 83
rect -28 77 -22 79
rect 12 79 14 81
rect 16 79 18 81
rect 85 81 91 83
rect 12 77 18 79
rect 85 79 87 81
rect 89 79 91 81
rect 116 81 122 83
rect 85 77 91 79
rect 116 79 118 81
rect 120 79 122 81
rect 189 81 195 83
rect 116 77 122 79
rect 189 79 191 81
rect 193 79 195 81
rect 257 81 263 83
rect 189 77 195 79
rect 257 79 259 81
rect 261 79 263 81
rect 305 81 311 83
rect 257 77 263 79
rect 305 79 307 81
rect 309 79 311 81
rect 305 77 311 79
<< nmos >>
rect -22 276 -20 285
rect -12 276 -10 282
rect -2 276 0 282
rect 18 278 20 287
rect 31 278 33 289
rect 38 278 40 289
rect 58 276 60 285
rect 74 281 76 290
rect 84 281 86 290
rect 94 281 96 293
rect 101 281 103 293
rect 122 278 124 287
rect 135 278 137 289
rect 142 278 144 289
rect 162 276 164 285
rect 178 281 180 290
rect 188 281 190 290
rect 198 281 200 293
rect 205 281 207 293
rect 235 278 237 289
rect 242 278 244 289
rect 255 278 257 287
rect 283 276 285 282
rect 293 276 295 282
rect 303 276 305 285
rect 332 281 334 290
rect 342 282 344 290
rect 349 282 351 290
rect 359 282 361 290
rect 366 282 368 290
rect 376 282 378 288
rect 406 281 408 290
rect 416 282 418 290
rect 423 282 425 290
rect 433 282 435 290
rect 440 282 442 290
rect 450 282 452 288
rect 480 281 482 290
rect 490 282 492 290
rect 497 282 499 290
rect 507 282 509 290
rect 514 282 516 290
rect 524 282 526 288
rect -22 175 -20 184
rect -12 178 -10 184
rect -2 178 0 184
rect 18 173 20 182
rect 31 171 33 182
rect 38 171 40 182
rect 58 175 60 184
rect 74 170 76 179
rect 84 170 86 179
rect 94 167 96 179
rect 101 167 103 179
rect 122 173 124 182
rect 135 171 137 182
rect 142 171 144 182
rect 162 175 164 184
rect 178 170 180 179
rect 188 170 190 179
rect 198 167 200 179
rect 205 167 207 179
rect 235 171 237 182
rect 242 171 244 182
rect 255 173 257 182
rect 283 178 285 184
rect 293 178 295 184
rect 303 175 305 184
rect 332 170 334 179
rect 342 170 344 178
rect 349 170 351 178
rect 359 170 361 178
rect 366 170 368 178
rect 376 172 378 178
rect 406 170 408 179
rect 416 170 418 178
rect 423 170 425 178
rect 433 170 435 178
rect 440 170 442 178
rect 450 172 452 178
rect 480 170 482 179
rect 490 170 492 178
rect 497 170 499 178
rect 507 170 509 178
rect 514 170 516 178
rect 524 172 526 178
rect -22 132 -20 141
rect -12 132 -10 138
rect -2 132 0 138
rect 18 134 20 143
rect 31 134 33 145
rect 38 134 40 145
rect 58 132 60 141
rect 74 137 76 146
rect 84 137 86 146
rect 94 137 96 149
rect 101 137 103 149
rect 122 134 124 143
rect 135 134 137 145
rect 142 134 144 145
rect 162 132 164 141
rect 178 137 180 146
rect 188 137 190 146
rect 198 137 200 149
rect 205 137 207 149
rect 235 134 237 145
rect 242 134 244 145
rect 255 134 257 143
rect 283 132 285 138
rect 293 132 295 138
rect 303 132 305 141
rect 332 137 334 146
rect 342 138 344 146
rect 349 138 351 146
rect 359 138 361 146
rect 366 138 368 146
rect 376 138 378 144
rect 406 137 408 146
rect 416 138 418 146
rect 423 138 425 146
rect 433 138 435 146
rect 440 138 442 146
rect 450 138 452 144
rect 480 137 482 146
rect 490 138 492 146
rect 497 138 499 146
rect 507 138 509 146
rect 514 138 516 146
rect 524 138 526 144
rect -22 31 -20 40
rect -12 34 -10 40
rect -2 34 0 40
rect 18 29 20 38
rect 31 27 33 38
rect 38 27 40 38
rect 58 31 60 40
rect 74 26 76 35
rect 84 26 86 35
rect 94 23 96 35
rect 101 23 103 35
rect 122 29 124 38
rect 135 27 137 38
rect 142 27 144 38
rect 162 31 164 40
rect 178 26 180 35
rect 188 26 190 35
rect 198 23 200 35
rect 205 23 207 35
rect 235 27 237 38
rect 242 27 244 38
rect 255 29 257 38
rect 283 34 285 40
rect 293 34 295 40
rect 303 31 305 40
rect 332 26 334 35
rect 342 26 344 34
rect 349 26 351 34
rect 359 26 361 34
rect 366 26 368 34
rect 376 28 378 34
rect 406 26 408 35
rect 416 26 418 34
rect 423 26 425 34
rect 433 26 435 34
rect 440 26 442 34
rect 450 28 452 34
rect 480 26 482 35
rect 490 26 492 34
rect 497 26 499 34
rect 507 26 509 34
rect 514 26 516 34
rect 524 28 526 34
<< pmos >>
rect -22 246 -20 264
rect -9 236 -7 257
rect -2 236 0 257
rect 18 245 20 263
rect 28 243 30 256
rect 38 243 40 256
rect 66 236 68 263
rect 82 245 84 263
rect 92 245 94 263
rect 102 236 104 263
rect 122 245 124 263
rect 132 243 134 256
rect 142 243 144 256
rect 170 236 172 263
rect 186 245 188 263
rect 196 245 198 263
rect 206 236 208 263
rect 235 243 237 256
rect 245 243 247 256
rect 255 245 257 263
rect 283 236 285 257
rect 290 236 292 257
rect 303 246 305 264
rect 332 236 334 254
rect 376 256 378 264
rect 342 236 344 252
rect 349 236 351 252
rect 359 236 361 252
rect 366 236 368 252
rect 406 236 408 254
rect 450 256 452 264
rect 416 236 418 252
rect 423 236 425 252
rect 433 236 435 252
rect 440 236 442 252
rect 480 236 482 254
rect 524 256 526 264
rect 490 236 492 252
rect 497 236 499 252
rect 507 236 509 252
rect 514 236 516 252
rect -22 196 -20 214
rect -9 203 -7 224
rect -2 203 0 224
rect 18 197 20 215
rect 28 204 30 217
rect 38 204 40 217
rect 66 197 68 224
rect 82 197 84 215
rect 92 197 94 215
rect 102 197 104 224
rect 122 197 124 215
rect 132 204 134 217
rect 142 204 144 217
rect 170 197 172 224
rect 186 197 188 215
rect 196 197 198 215
rect 206 197 208 224
rect 235 204 237 217
rect 245 204 247 217
rect 255 197 257 215
rect 283 203 285 224
rect 290 203 292 224
rect 303 196 305 214
rect 332 206 334 224
rect 342 208 344 224
rect 349 208 351 224
rect 359 208 361 224
rect 366 208 368 224
rect 406 206 408 224
rect 416 208 418 224
rect 423 208 425 224
rect 433 208 435 224
rect 440 208 442 224
rect 376 196 378 204
rect 480 206 482 224
rect 490 208 492 224
rect 497 208 499 224
rect 507 208 509 224
rect 514 208 516 224
rect 450 196 452 204
rect 524 196 526 204
rect -22 102 -20 120
rect -9 92 -7 113
rect -2 92 0 113
rect 18 101 20 119
rect 28 99 30 112
rect 38 99 40 112
rect 66 92 68 119
rect 82 101 84 119
rect 92 101 94 119
rect 102 92 104 119
rect 122 101 124 119
rect 132 99 134 112
rect 142 99 144 112
rect 170 92 172 119
rect 186 101 188 119
rect 196 101 198 119
rect 206 92 208 119
rect 235 99 237 112
rect 245 99 247 112
rect 255 101 257 119
rect 283 92 285 113
rect 290 92 292 113
rect 303 102 305 120
rect 332 92 334 110
rect 376 112 378 120
rect 342 92 344 108
rect 349 92 351 108
rect 359 92 361 108
rect 366 92 368 108
rect 406 92 408 110
rect 450 112 452 120
rect 416 92 418 108
rect 423 92 425 108
rect 433 92 435 108
rect 440 92 442 108
rect 480 92 482 110
rect 524 112 526 120
rect 490 92 492 108
rect 497 92 499 108
rect 507 92 509 108
rect 514 92 516 108
rect -22 52 -20 70
rect -9 59 -7 80
rect -2 59 0 80
rect 18 53 20 71
rect 28 60 30 73
rect 38 60 40 73
rect 66 53 68 80
rect 82 53 84 71
rect 92 53 94 71
rect 102 53 104 80
rect 122 53 124 71
rect 132 60 134 73
rect 142 60 144 73
rect 170 53 172 80
rect 186 53 188 71
rect 196 53 198 71
rect 206 53 208 80
rect 235 60 237 73
rect 245 60 247 73
rect 255 53 257 71
rect 283 59 285 80
rect 290 59 292 80
rect 303 52 305 70
rect 332 62 334 80
rect 342 64 344 80
rect 349 64 351 80
rect 359 64 361 80
rect 366 64 368 80
rect 406 62 408 80
rect 416 64 418 80
rect 423 64 425 80
rect 433 64 435 80
rect 440 64 442 80
rect 376 52 378 60
rect 480 62 482 80
rect 490 64 492 80
rect 497 64 499 80
rect 507 64 509 80
rect 514 64 516 80
rect 450 52 452 60
rect 524 52 526 60
<< polyct0 >>
rect -20 269 -18 271
rect 20 269 22 271
rect 90 269 92 271
rect 100 268 102 270
rect 124 269 126 271
rect 194 269 196 271
rect 204 268 206 270
rect 253 269 255 271
rect 333 274 335 276
rect 301 269 303 271
rect 351 275 353 277
rect 358 259 360 261
rect 407 274 409 276
rect 425 275 427 277
rect 432 259 434 261
rect 481 274 483 276
rect 499 275 501 277
rect 506 259 508 261
rect -20 189 -18 191
rect 20 189 22 191
rect 90 189 92 191
rect 100 190 102 192
rect 124 189 126 191
rect 194 189 196 191
rect 204 190 206 192
rect 253 189 255 191
rect 301 189 303 191
rect 358 199 360 201
rect 333 184 335 186
rect 351 183 353 185
rect 432 199 434 201
rect 407 184 409 186
rect 425 183 427 185
rect 506 199 508 201
rect 481 184 483 186
rect 499 183 501 185
rect -20 125 -18 127
rect 20 125 22 127
rect 90 125 92 127
rect 100 124 102 126
rect 124 125 126 127
rect 194 125 196 127
rect 204 124 206 126
rect 253 125 255 127
rect 333 130 335 132
rect 301 125 303 127
rect 351 131 353 133
rect 358 115 360 117
rect 407 130 409 132
rect 425 131 427 133
rect 432 115 434 117
rect 481 130 483 132
rect 499 131 501 133
rect 506 115 508 117
rect -20 45 -18 47
rect 20 45 22 47
rect 90 45 92 47
rect 100 46 102 48
rect 124 45 126 47
rect 194 45 196 47
rect 204 46 206 48
rect 253 45 255 47
rect 301 45 303 47
rect 358 55 360 57
rect 333 40 335 42
rect 351 39 353 41
rect 432 55 434 57
rect 407 40 409 42
rect 425 39 427 41
rect 506 55 508 57
rect 481 40 483 42
rect 499 39 501 41
<< polyct1 >>
rect -10 269 -8 271
rect 30 269 32 271
rect 0 262 2 264
rect 69 274 71 276
rect 40 261 42 263
rect 134 269 136 271
rect 53 261 55 263
rect 173 274 175 276
rect 144 261 146 263
rect 243 269 245 271
rect 157 261 159 263
rect 233 261 235 263
rect 291 269 293 271
rect 281 262 283 264
rect 341 264 343 266
rect 368 274 370 276
rect 415 264 417 266
rect 442 269 444 271
rect 381 249 383 251
rect 489 264 491 266
rect 516 269 518 271
rect 455 249 457 251
rect 529 249 531 251
rect 0 196 2 198
rect -10 189 -8 191
rect 40 197 42 199
rect 53 197 55 199
rect 30 189 32 191
rect 144 197 146 199
rect 157 197 159 199
rect 233 197 235 199
rect 69 184 71 186
rect 134 189 136 191
rect 173 184 175 186
rect 281 196 283 198
rect 243 189 245 191
rect 381 209 383 211
rect 291 189 293 191
rect 341 194 343 196
rect 455 209 457 211
rect 368 184 370 186
rect 415 194 417 196
rect 529 209 531 211
rect 442 189 444 191
rect 489 194 491 196
rect 516 189 518 191
rect -10 125 -8 127
rect 30 125 32 127
rect 0 118 2 120
rect 69 130 71 132
rect 40 117 42 119
rect 134 125 136 127
rect 53 117 55 119
rect 173 130 175 132
rect 144 117 146 119
rect 243 125 245 127
rect 157 117 159 119
rect 233 117 235 119
rect 291 125 293 127
rect 281 118 283 120
rect 341 120 343 122
rect 368 130 370 132
rect 415 120 417 122
rect 442 125 444 127
rect 381 105 383 107
rect 489 120 491 122
rect 516 125 518 127
rect 455 105 457 107
rect 529 105 531 107
rect 0 52 2 54
rect -10 45 -8 47
rect 40 53 42 55
rect 53 53 55 55
rect 30 45 32 47
rect 144 53 146 55
rect 157 53 159 55
rect 233 53 235 55
rect 69 40 71 42
rect 134 45 136 47
rect 173 40 175 42
rect 281 52 283 54
rect 243 45 245 47
rect 381 65 383 67
rect 291 45 293 47
rect 341 50 343 52
rect 455 65 457 67
rect 368 40 370 42
rect 415 50 417 52
rect 529 65 531 67
rect 442 45 444 47
rect 489 50 491 52
rect 516 45 518 47
<< ndifct0 >>
rect -16 291 -14 293
rect 3 291 5 293
rect -7 278 -5 280
rect 43 285 45 287
rect 67 286 69 288
rect 53 278 55 280
rect 79 283 81 285
rect 147 285 149 287
rect 171 286 173 288
rect 157 278 159 280
rect 183 283 185 285
rect 278 291 280 293
rect 230 285 232 287
rect 297 291 299 293
rect 288 278 290 280
rect 337 286 339 288
rect 354 286 356 288
rect 371 284 373 286
rect 381 284 383 286
rect 411 286 413 288
rect 428 286 430 288
rect 445 284 447 286
rect 455 284 457 286
rect 485 286 487 288
rect 502 286 504 288
rect 519 284 521 286
rect 529 284 531 286
rect -7 180 -5 182
rect -16 167 -14 169
rect 53 180 55 182
rect 43 173 45 175
rect 67 172 69 174
rect 3 167 5 169
rect 79 175 81 177
rect 157 180 159 182
rect 147 173 149 175
rect 171 172 173 174
rect 183 175 185 177
rect 230 173 232 175
rect 288 180 290 182
rect 278 167 280 169
rect 337 172 339 174
rect 354 172 356 174
rect 371 174 373 176
rect 381 174 383 176
rect 297 167 299 169
rect 411 172 413 174
rect 428 172 430 174
rect 445 174 447 176
rect 455 174 457 176
rect 485 172 487 174
rect 502 172 504 174
rect 519 174 521 176
rect 529 174 531 176
rect -16 147 -14 149
rect 3 147 5 149
rect -7 134 -5 136
rect 43 141 45 143
rect 67 142 69 144
rect 53 134 55 136
rect 79 139 81 141
rect 147 141 149 143
rect 171 142 173 144
rect 157 134 159 136
rect 183 139 185 141
rect 278 147 280 149
rect 230 141 232 143
rect 297 147 299 149
rect 288 134 290 136
rect 337 142 339 144
rect 354 142 356 144
rect 371 140 373 142
rect 381 140 383 142
rect 411 142 413 144
rect 428 142 430 144
rect 445 140 447 142
rect 455 140 457 142
rect 485 142 487 144
rect 502 142 504 144
rect 519 140 521 142
rect 529 140 531 142
rect -7 36 -5 38
rect -16 23 -14 25
rect 53 36 55 38
rect 43 29 45 31
rect 67 28 69 30
rect 3 23 5 25
rect 79 31 81 33
rect 157 36 159 38
rect 147 29 149 31
rect 171 28 173 30
rect 183 31 185 33
rect 230 29 232 31
rect 288 36 290 38
rect 278 23 280 25
rect 337 28 339 30
rect 354 28 356 30
rect 371 30 373 32
rect 381 30 383 32
rect 297 23 299 25
rect 411 28 413 30
rect 428 28 430 30
rect 445 30 447 32
rect 455 30 457 32
rect 485 28 487 30
rect 502 28 504 30
rect 519 30 521 32
rect 529 30 531 32
<< ndifct1 >>
rect 24 295 26 297
rect -27 278 -25 280
rect 107 295 109 297
rect 128 295 130 297
rect 13 283 15 285
rect 89 285 91 287
rect 211 295 213 297
rect 249 295 251 297
rect 117 283 119 285
rect 193 285 195 287
rect 260 283 262 285
rect 327 283 329 285
rect 401 283 403 285
rect 308 278 310 280
rect 475 283 477 285
rect -27 180 -25 182
rect 13 175 15 177
rect 89 173 91 175
rect 24 163 26 165
rect 117 175 119 177
rect 107 163 109 165
rect 193 173 195 175
rect 128 163 130 165
rect 260 175 262 177
rect 211 163 213 165
rect 308 180 310 182
rect 327 175 329 177
rect 249 163 251 165
rect 401 175 403 177
rect 475 175 477 177
rect 24 151 26 153
rect -27 134 -25 136
rect 107 151 109 153
rect 128 151 130 153
rect 13 139 15 141
rect 89 141 91 143
rect 211 151 213 153
rect 249 151 251 153
rect 117 139 119 141
rect 193 141 195 143
rect 260 139 262 141
rect 327 139 329 141
rect 401 139 403 141
rect 308 134 310 136
rect 475 139 477 141
rect -27 36 -25 38
rect 13 31 15 33
rect 89 29 91 31
rect 24 19 26 21
rect 117 31 119 33
rect 107 19 109 21
rect 193 29 195 31
rect 128 19 130 21
rect 260 31 262 33
rect 211 19 213 21
rect 308 36 310 38
rect 327 31 329 33
rect 249 19 251 21
rect 401 31 403 33
rect 475 31 477 33
<< ntiect1 >>
rect -26 235 -24 237
rect 14 235 16 237
rect 87 235 89 237
rect 118 235 120 237
rect 191 235 193 237
rect 259 235 261 237
rect 307 235 309 237
rect -26 223 -24 225
rect 14 223 16 225
rect 87 223 89 225
rect 118 223 120 225
rect 191 223 193 225
rect 259 223 261 225
rect 307 223 309 225
rect -26 91 -24 93
rect 14 91 16 93
rect 87 91 89 93
rect 118 91 120 93
rect 191 91 193 93
rect 259 91 261 93
rect 307 91 309 93
rect -26 79 -24 81
rect 14 79 16 81
rect 87 79 89 81
rect 118 79 120 81
rect 191 79 193 81
rect 259 79 261 81
rect 307 79 309 81
<< ptiect1 >>
rect -26 295 -24 297
rect 14 295 16 297
rect 54 295 56 297
rect 118 295 120 297
rect 158 295 160 297
rect 259 295 261 297
rect 307 295 309 297
rect -26 163 -24 165
rect 14 163 16 165
rect 54 163 56 165
rect 118 163 120 165
rect 158 163 160 165
rect 259 163 261 165
rect 307 163 309 165
rect -26 151 -24 153
rect 14 151 16 153
rect 54 151 56 153
rect 118 151 120 153
rect 158 151 160 153
rect 259 151 261 153
rect 307 151 309 153
rect -26 19 -24 21
rect 14 19 16 21
rect 54 19 56 21
rect 118 19 120 21
rect 158 19 160 21
rect 259 19 261 21
rect 307 19 309 21
<< pdifct0 >>
rect -16 238 -14 240
rect 3 245 5 247
rect 61 259 63 261
rect 23 247 25 249
rect 33 252 35 254
rect 33 245 35 247
rect 43 245 45 247
rect 71 245 73 247
rect 87 259 89 261
rect 87 252 89 254
rect 71 238 73 240
rect 107 244 109 246
rect 165 259 167 261
rect 127 247 129 249
rect 137 252 139 254
rect 137 245 139 247
rect 147 245 149 247
rect 175 245 177 247
rect 191 259 193 261
rect 191 252 193 254
rect 175 238 177 240
rect 211 244 213 246
rect 230 245 232 247
rect 240 252 242 254
rect 240 245 242 247
rect 250 247 252 249
rect 278 245 280 247
rect 297 238 299 240
rect 381 260 383 262
rect 337 238 339 240
rect 354 248 356 250
rect 371 238 373 240
rect 455 260 457 262
rect 411 238 413 240
rect 428 248 430 250
rect 445 238 447 240
rect 529 260 531 262
rect 485 238 487 240
rect 502 248 504 250
rect 519 238 521 240
rect -16 220 -14 222
rect 3 213 5 215
rect 23 211 25 213
rect 33 213 35 215
rect 33 206 35 208
rect 43 213 45 215
rect 61 199 63 201
rect 71 220 73 222
rect 71 213 73 215
rect 87 206 89 208
rect 87 199 89 201
rect 107 214 109 216
rect 127 211 129 213
rect 137 213 139 215
rect 137 206 139 208
rect 147 213 149 215
rect 165 199 167 201
rect 175 220 177 222
rect 175 213 177 215
rect 191 206 193 208
rect 191 199 193 201
rect 211 214 213 216
rect 230 213 232 215
rect 240 213 242 215
rect 240 206 242 208
rect 250 211 252 213
rect 278 213 280 215
rect 297 220 299 222
rect 337 220 339 222
rect 354 210 356 212
rect 371 220 373 222
rect 411 220 413 222
rect 428 210 430 212
rect 445 220 447 222
rect 381 198 383 200
rect 485 220 487 222
rect 502 210 504 212
rect 519 220 521 222
rect 455 198 457 200
rect 529 198 531 200
rect -16 94 -14 96
rect 3 101 5 103
rect 61 115 63 117
rect 23 103 25 105
rect 33 108 35 110
rect 33 101 35 103
rect 43 101 45 103
rect 71 101 73 103
rect 87 115 89 117
rect 87 108 89 110
rect 71 94 73 96
rect 107 100 109 102
rect 165 115 167 117
rect 127 103 129 105
rect 137 108 139 110
rect 137 101 139 103
rect 147 101 149 103
rect 175 101 177 103
rect 191 115 193 117
rect 191 108 193 110
rect 175 94 177 96
rect 211 100 213 102
rect 230 101 232 103
rect 240 108 242 110
rect 240 101 242 103
rect 250 103 252 105
rect 278 101 280 103
rect 297 94 299 96
rect 381 116 383 118
rect 337 94 339 96
rect 354 104 356 106
rect 371 94 373 96
rect 455 116 457 118
rect 411 94 413 96
rect 428 104 430 106
rect 445 94 447 96
rect 529 116 531 118
rect 485 94 487 96
rect 502 104 504 106
rect 519 94 521 96
rect -16 76 -14 78
rect 3 69 5 71
rect 23 67 25 69
rect 33 69 35 71
rect 33 62 35 64
rect 43 69 45 71
rect 61 55 63 57
rect 71 76 73 78
rect 71 69 73 71
rect 87 62 89 64
rect 87 55 89 57
rect 107 70 109 72
rect 127 67 129 69
rect 137 69 139 71
rect 137 62 139 64
rect 147 69 149 71
rect 165 55 167 57
rect 175 76 177 78
rect 175 69 177 71
rect 191 62 193 64
rect 191 55 193 57
rect 211 70 213 72
rect 230 69 232 71
rect 240 69 242 71
rect 240 62 242 64
rect 250 67 252 69
rect 278 69 280 71
rect 297 76 299 78
rect 337 76 339 78
rect 354 66 356 68
rect 371 76 373 78
rect 411 76 413 78
rect 428 66 430 68
rect 445 76 447 78
rect 381 54 383 56
rect 485 76 487 78
rect 502 66 504 68
rect 519 76 521 78
rect 455 54 457 56
rect 529 54 531 56
<< pdifct1 >>
rect -27 255 -25 257
rect -27 248 -25 250
rect 13 259 15 261
rect 13 252 15 254
rect 97 252 99 254
rect 117 259 119 261
rect 117 252 119 254
rect 201 252 203 254
rect 260 259 262 261
rect 260 252 262 254
rect 308 255 310 257
rect 308 248 310 250
rect 327 245 329 247
rect 401 245 403 247
rect 475 245 477 247
rect -27 210 -25 212
rect -27 203 -25 205
rect 13 206 15 208
rect 13 199 15 201
rect 97 206 99 208
rect 117 206 119 208
rect 117 199 119 201
rect 201 206 203 208
rect 260 206 262 208
rect 260 199 262 201
rect 308 210 310 212
rect 327 213 329 215
rect 401 213 403 215
rect 308 203 310 205
rect 475 213 477 215
rect -27 111 -25 113
rect -27 104 -25 106
rect 13 115 15 117
rect 13 108 15 110
rect 97 108 99 110
rect 117 115 119 117
rect 117 108 119 110
rect 201 108 203 110
rect 260 115 262 117
rect 260 108 262 110
rect 308 111 310 113
rect 308 104 310 106
rect 327 101 329 103
rect 401 101 403 103
rect 475 101 477 103
rect -27 66 -25 68
rect -27 59 -25 61
rect 13 62 15 64
rect 13 55 15 57
rect 97 62 99 64
rect 117 62 119 64
rect 117 55 119 57
rect 201 62 203 64
rect 260 62 262 64
rect 260 55 262 57
rect 308 66 310 68
rect 327 69 329 71
rect 401 69 403 71
rect 308 59 310 61
rect 475 69 477 71
<< alu0 >>
rect -18 293 -12 294
rect -18 291 -16 293
rect -14 291 -12 293
rect -18 290 -12 291
rect 1 293 7 294
rect 1 291 3 293
rect 5 291 7 293
rect 1 290 7 291
rect 65 288 71 294
rect 27 287 47 288
rect 27 285 43 287
rect 45 285 47 287
rect 65 286 67 288
rect 69 286 71 288
rect 65 285 71 286
rect 78 285 82 287
rect 27 284 47 285
rect -21 280 -3 281
rect -21 278 -7 280
rect -5 278 -3 280
rect -21 277 -3 278
rect -21 271 -17 277
rect -21 269 -20 271
rect -18 269 -17 271
rect -25 248 -24 259
rect -21 256 -17 269
rect -2 264 4 265
rect -21 252 -6 256
rect -10 248 -6 252
rect 15 281 16 283
rect 27 280 31 284
rect 78 283 79 285
rect 81 283 82 285
rect 19 276 31 280
rect 19 271 23 276
rect 19 269 20 271
rect 22 269 23 271
rect 19 257 23 269
rect 52 280 56 282
rect 52 278 53 280
rect 55 278 56 280
rect 52 272 56 278
rect 78 280 82 283
rect 78 276 102 280
rect 52 268 63 272
rect 19 254 36 257
rect 19 253 33 254
rect 32 252 33 253
rect 35 252 36 254
rect 21 249 27 250
rect -10 247 7 248
rect -10 245 3 247
rect 5 245 7 247
rect -10 244 7 245
rect 21 247 23 249
rect 25 247 27 249
rect -18 240 -12 241
rect -18 238 -16 240
rect -14 238 -12 240
rect 21 238 27 247
rect 32 247 36 252
rect 59 262 63 268
rect 98 272 102 276
rect 78 271 94 272
rect 78 269 90 271
rect 92 269 94 271
rect 78 268 94 269
rect 98 270 103 272
rect 98 268 100 270
rect 102 268 103 270
rect 78 262 82 268
rect 98 266 103 268
rect 98 264 102 266
rect 59 261 82 262
rect 59 259 61 261
rect 63 259 82 261
rect 59 258 82 259
rect 32 245 33 247
rect 35 245 36 247
rect 32 243 36 245
rect 41 247 47 248
rect 41 245 43 247
rect 45 245 47 247
rect 41 238 47 245
rect 70 247 74 249
rect 70 245 71 247
rect 73 245 74 247
rect 70 240 74 245
rect 78 247 82 258
rect 86 261 102 264
rect 86 259 87 261
rect 89 260 102 261
rect 89 259 90 260
rect 86 254 90 259
rect 86 252 87 254
rect 89 252 90 254
rect 86 250 90 252
rect 169 288 175 294
rect 276 293 282 294
rect 276 291 278 293
rect 280 291 282 293
rect 276 290 282 291
rect 295 293 301 294
rect 295 291 297 293
rect 299 291 301 293
rect 295 290 301 291
rect 131 287 151 288
rect 131 285 147 287
rect 149 285 151 287
rect 169 286 171 288
rect 173 286 175 288
rect 169 285 175 286
rect 182 285 186 287
rect 131 284 151 285
rect 119 281 120 283
rect 131 280 135 284
rect 182 283 183 285
rect 185 283 186 285
rect 228 287 248 288
rect 228 285 230 287
rect 232 285 248 287
rect 228 284 248 285
rect 123 276 135 280
rect 123 271 127 276
rect 123 269 124 271
rect 126 269 127 271
rect 123 257 127 269
rect 156 280 160 282
rect 156 278 157 280
rect 159 278 160 280
rect 156 272 160 278
rect 182 280 186 283
rect 182 276 206 280
rect 156 268 167 272
rect 123 254 140 257
rect 123 253 137 254
rect 136 252 137 253
rect 139 252 140 254
rect 125 249 131 250
rect 125 247 127 249
rect 129 247 131 249
rect 78 246 111 247
rect 78 244 107 246
rect 109 244 111 246
rect 78 243 111 244
rect 70 238 71 240
rect 73 238 74 240
rect 125 238 131 247
rect 136 247 140 252
rect 163 262 167 268
rect 202 272 206 276
rect 182 271 198 272
rect 182 269 194 271
rect 196 269 198 271
rect 182 268 198 269
rect 202 270 207 272
rect 202 268 204 270
rect 206 268 207 270
rect 182 262 186 268
rect 202 266 207 268
rect 202 264 206 266
rect 163 261 186 262
rect 163 259 165 261
rect 167 259 186 261
rect 163 258 186 259
rect 136 245 137 247
rect 139 245 140 247
rect 136 243 140 245
rect 145 247 151 248
rect 145 245 147 247
rect 149 245 151 247
rect 145 238 151 245
rect 174 247 178 249
rect 174 245 175 247
rect 177 245 178 247
rect 174 240 178 245
rect 182 247 186 258
rect 190 261 206 264
rect 190 259 191 261
rect 193 260 206 261
rect 193 259 194 260
rect 190 254 194 259
rect 244 280 248 284
rect 259 281 260 283
rect 244 276 256 280
rect 252 271 256 276
rect 252 269 253 271
rect 255 269 256 271
rect 190 252 191 254
rect 193 252 194 254
rect 190 250 194 252
rect 252 257 256 269
rect 336 288 340 294
rect 336 286 337 288
rect 339 286 340 288
rect 336 284 340 286
rect 343 288 358 289
rect 343 286 354 288
rect 356 286 358 288
rect 343 285 358 286
rect 369 286 375 294
rect 410 288 414 294
rect 286 280 304 281
rect 286 278 288 280
rect 290 278 304 280
rect 286 277 304 278
rect 300 271 304 277
rect 300 269 301 271
rect 303 269 304 271
rect 279 264 285 265
rect 239 254 256 257
rect 239 252 240 254
rect 242 253 256 254
rect 242 252 243 253
rect 228 247 234 248
rect 182 246 215 247
rect 182 244 211 246
rect 213 244 215 246
rect 182 243 215 244
rect 228 245 230 247
rect 232 245 234 247
rect 174 238 175 240
rect 177 238 178 240
rect 228 238 234 245
rect 239 247 243 252
rect 300 256 304 269
rect 289 252 304 256
rect 239 245 240 247
rect 242 245 243 247
rect 239 243 243 245
rect 248 249 254 250
rect 248 247 250 249
rect 252 247 254 249
rect 289 248 293 252
rect 307 248 308 259
rect 248 238 254 247
rect 276 247 293 248
rect 276 245 278 247
rect 280 245 293 247
rect 276 244 293 245
rect 343 280 347 285
rect 369 284 371 286
rect 373 284 375 286
rect 369 283 375 284
rect 379 286 385 287
rect 379 284 381 286
rect 383 284 385 286
rect 379 283 385 284
rect 333 278 347 280
rect 332 276 347 278
rect 350 277 361 279
rect 332 274 333 276
rect 335 274 337 276
rect 332 272 337 274
rect 350 275 351 277
rect 353 275 361 277
rect 350 273 361 275
rect 333 267 337 272
rect 333 265 334 267
rect 336 265 337 267
rect 333 255 337 265
rect 357 263 361 273
rect 381 263 385 283
rect 357 262 385 263
rect 357 261 370 262
rect 357 259 358 261
rect 360 260 370 261
rect 372 260 381 262
rect 383 260 385 262
rect 360 259 385 260
rect 410 286 411 288
rect 413 286 414 288
rect 410 284 414 286
rect 417 288 432 289
rect 417 286 428 288
rect 430 286 432 288
rect 417 285 432 286
rect 443 286 449 294
rect 484 288 488 294
rect 417 280 421 285
rect 443 284 445 286
rect 447 284 449 286
rect 443 283 449 284
rect 453 286 459 287
rect 453 284 455 286
rect 457 284 459 286
rect 453 283 459 284
rect 407 278 421 280
rect 406 276 421 278
rect 424 277 435 279
rect 406 274 407 276
rect 409 274 411 276
rect 406 272 411 274
rect 424 275 425 277
rect 427 275 435 277
rect 424 273 435 275
rect 357 257 361 259
rect 333 251 349 255
rect 345 250 358 251
rect 345 248 354 250
rect 356 248 358 250
rect 345 247 358 248
rect 407 267 411 272
rect 407 265 408 267
rect 410 265 411 267
rect 407 255 411 265
rect 431 263 435 273
rect 455 263 459 283
rect 431 262 459 263
rect 431 261 444 262
rect 431 259 432 261
rect 434 260 444 261
rect 446 260 455 262
rect 457 260 459 262
rect 434 259 459 260
rect 484 286 485 288
rect 487 286 488 288
rect 484 284 488 286
rect 491 288 506 289
rect 491 286 502 288
rect 504 286 506 288
rect 491 285 506 286
rect 517 286 523 294
rect 431 257 435 259
rect 407 251 423 255
rect 419 250 432 251
rect 419 248 428 250
rect 430 248 432 250
rect 419 247 432 248
rect 491 280 495 285
rect 517 284 519 286
rect 521 284 523 286
rect 517 283 523 284
rect 527 286 533 287
rect 527 284 529 286
rect 531 284 533 286
rect 527 283 533 284
rect 481 278 495 280
rect 480 276 495 278
rect 498 277 509 279
rect 480 274 481 276
rect 483 274 485 276
rect 480 272 485 274
rect 498 275 499 277
rect 501 275 509 277
rect 498 273 509 275
rect 481 267 485 272
rect 481 265 482 267
rect 484 265 485 267
rect 481 255 485 265
rect 488 262 489 268
rect 505 263 509 273
rect 529 263 533 283
rect 505 262 533 263
rect 505 261 518 262
rect 505 259 506 261
rect 508 260 518 261
rect 520 260 529 262
rect 531 260 533 262
rect 508 259 533 260
rect 505 257 509 259
rect 481 251 497 255
rect 493 250 506 251
rect 493 248 502 250
rect 504 248 506 250
rect 493 247 506 248
rect 295 240 301 241
rect 295 238 297 240
rect 299 238 301 240
rect 335 240 341 241
rect 335 238 337 240
rect 339 238 341 240
rect 370 240 374 242
rect 370 238 371 240
rect 373 238 374 240
rect 409 240 415 241
rect 409 238 411 240
rect 413 238 415 240
rect 444 240 448 242
rect 444 238 445 240
rect 447 238 448 240
rect 483 240 489 241
rect 483 238 485 240
rect 487 238 489 240
rect 518 240 522 242
rect 518 238 519 240
rect 521 238 522 240
rect -18 220 -16 222
rect -14 220 -12 222
rect -18 219 -12 220
rect -10 215 7 216
rect -10 213 3 215
rect 5 213 7 215
rect -10 212 7 213
rect 21 213 27 222
rect -25 201 -24 212
rect -10 208 -6 212
rect 21 211 23 213
rect 25 211 27 213
rect 21 210 27 211
rect 32 215 36 217
rect 32 213 33 215
rect 35 213 36 215
rect -21 204 -6 208
rect -21 191 -17 204
rect 32 208 36 213
rect 41 215 47 222
rect 70 220 71 222
rect 73 220 74 222
rect 41 213 43 215
rect 45 213 47 215
rect 41 212 47 213
rect 70 215 74 220
rect 70 213 71 215
rect 73 213 74 215
rect 70 211 74 213
rect 78 216 111 217
rect 78 214 107 216
rect 109 214 111 216
rect 78 213 111 214
rect 125 213 131 222
rect 32 207 33 208
rect 19 206 33 207
rect 35 206 36 208
rect 19 203 36 206
rect -2 195 4 196
rect -21 189 -20 191
rect -18 189 -17 191
rect -21 183 -17 189
rect -21 182 -3 183
rect -21 180 -7 182
rect -5 180 -3 182
rect -21 179 -3 180
rect 19 191 23 203
rect 78 202 82 213
rect 125 211 127 213
rect 129 211 131 213
rect 125 210 131 211
rect 136 215 140 217
rect 136 213 137 215
rect 139 213 140 215
rect 59 201 82 202
rect 59 199 61 201
rect 63 199 82 201
rect 59 198 82 199
rect 59 192 63 198
rect 19 189 20 191
rect 22 189 23 191
rect 19 184 23 189
rect 19 180 31 184
rect 15 177 16 179
rect 27 176 31 180
rect 52 188 63 192
rect 52 182 56 188
rect 78 192 82 198
rect 86 208 90 210
rect 86 206 87 208
rect 89 206 90 208
rect 86 201 90 206
rect 86 199 87 201
rect 89 200 90 201
rect 89 199 102 200
rect 86 196 102 199
rect 98 194 102 196
rect 98 192 103 194
rect 78 191 94 192
rect 78 189 90 191
rect 92 189 94 191
rect 78 188 94 189
rect 98 190 100 192
rect 102 190 103 192
rect 98 188 103 190
rect 52 180 53 182
rect 55 180 56 182
rect 52 178 56 180
rect 98 184 102 188
rect 78 180 102 184
rect 78 177 82 180
rect 27 175 47 176
rect 78 175 79 177
rect 81 175 82 177
rect 27 173 43 175
rect 45 173 47 175
rect 27 172 47 173
rect 65 174 71 175
rect 65 172 67 174
rect 69 172 71 174
rect 78 173 82 175
rect 136 208 140 213
rect 145 215 151 222
rect 174 220 175 222
rect 177 220 178 222
rect 145 213 147 215
rect 149 213 151 215
rect 145 212 151 213
rect 174 215 178 220
rect 174 213 175 215
rect 177 213 178 215
rect 174 211 178 213
rect 182 216 215 217
rect 182 214 211 216
rect 213 214 215 216
rect 182 213 215 214
rect 228 215 234 222
rect 228 213 230 215
rect 232 213 234 215
rect 136 207 137 208
rect 123 206 137 207
rect 139 206 140 208
rect 123 203 140 206
rect 123 191 127 203
rect 182 202 186 213
rect 228 212 234 213
rect 239 215 243 217
rect 239 213 240 215
rect 242 213 243 215
rect 163 201 186 202
rect 163 199 165 201
rect 167 199 186 201
rect 163 198 186 199
rect 163 192 167 198
rect 123 189 124 191
rect 126 189 127 191
rect 123 184 127 189
rect 123 180 135 184
rect 119 177 120 179
rect -18 169 -12 170
rect -18 167 -16 169
rect -14 167 -12 169
rect -18 166 -12 167
rect 1 169 7 170
rect 1 167 3 169
rect 5 167 7 169
rect 1 166 7 167
rect 65 166 71 172
rect 131 176 135 180
rect 156 188 167 192
rect 156 182 160 188
rect 182 192 186 198
rect 190 208 194 210
rect 190 206 191 208
rect 193 206 194 208
rect 190 201 194 206
rect 190 199 191 201
rect 193 200 194 201
rect 193 199 206 200
rect 190 196 206 199
rect 202 194 206 196
rect 202 192 207 194
rect 182 191 198 192
rect 182 189 194 191
rect 196 189 198 191
rect 182 188 198 189
rect 202 190 204 192
rect 206 190 207 192
rect 202 188 207 190
rect 156 180 157 182
rect 159 180 160 182
rect 156 178 160 180
rect 202 184 206 188
rect 182 180 206 184
rect 239 208 243 213
rect 248 213 254 222
rect 295 220 297 222
rect 299 220 301 222
rect 295 219 301 220
rect 335 220 337 222
rect 339 220 341 222
rect 335 219 341 220
rect 370 220 371 222
rect 373 220 374 222
rect 370 218 374 220
rect 409 220 411 222
rect 413 220 415 222
rect 409 219 415 220
rect 444 220 445 222
rect 447 220 448 222
rect 444 218 448 220
rect 483 220 485 222
rect 487 220 489 222
rect 483 219 489 220
rect 518 220 519 222
rect 521 220 522 222
rect 518 218 522 220
rect 248 211 250 213
rect 252 211 254 213
rect 276 215 293 216
rect 276 213 278 215
rect 280 213 293 215
rect 276 212 293 213
rect 248 210 254 211
rect 239 206 240 208
rect 242 207 243 208
rect 242 206 256 207
rect 239 203 256 206
rect 182 177 186 180
rect 131 175 151 176
rect 182 175 183 177
rect 185 175 186 177
rect 252 191 256 203
rect 252 189 253 191
rect 255 189 256 191
rect 252 184 256 189
rect 244 180 256 184
rect 289 208 293 212
rect 289 204 304 208
rect 279 195 285 196
rect 244 176 248 180
rect 259 177 260 179
rect 300 191 304 204
rect 307 201 308 212
rect 300 189 301 191
rect 303 189 304 191
rect 300 183 304 189
rect 286 182 304 183
rect 286 180 288 182
rect 290 180 304 182
rect 286 179 304 180
rect 345 212 358 213
rect 345 210 354 212
rect 356 210 358 212
rect 345 209 358 210
rect 333 205 349 209
rect 333 195 337 205
rect 419 212 432 213
rect 357 201 361 203
rect 333 193 334 195
rect 336 193 337 195
rect 333 188 337 193
rect 332 186 337 188
rect 357 199 358 201
rect 360 200 385 201
rect 360 199 370 200
rect 357 198 370 199
rect 372 198 381 200
rect 383 198 385 200
rect 357 197 385 198
rect 357 187 361 197
rect 332 184 333 186
rect 335 184 337 186
rect 350 185 361 187
rect 332 182 347 184
rect 333 180 347 182
rect 350 183 351 185
rect 353 183 361 185
rect 350 181 361 183
rect 131 173 147 175
rect 149 173 151 175
rect 131 172 151 173
rect 169 174 175 175
rect 169 172 171 174
rect 173 172 175 174
rect 182 173 186 175
rect 228 175 248 176
rect 228 173 230 175
rect 232 173 248 175
rect 228 172 248 173
rect 169 166 175 172
rect 336 174 340 176
rect 336 172 337 174
rect 339 172 340 174
rect 276 169 282 170
rect 276 167 278 169
rect 280 167 282 169
rect 276 166 282 167
rect 295 169 301 170
rect 295 167 297 169
rect 299 167 301 169
rect 295 166 301 167
rect 336 166 340 172
rect 343 175 347 180
rect 381 177 385 197
rect 369 176 375 177
rect 343 174 358 175
rect 343 172 354 174
rect 356 172 358 174
rect 343 171 358 172
rect 369 174 371 176
rect 373 174 375 176
rect 369 166 375 174
rect 379 176 385 177
rect 379 174 381 176
rect 383 174 385 176
rect 379 173 385 174
rect 419 210 428 212
rect 430 210 432 212
rect 419 209 432 210
rect 407 205 423 209
rect 407 195 411 205
rect 493 212 506 213
rect 431 201 435 203
rect 407 193 408 195
rect 410 193 411 195
rect 407 188 411 193
rect 431 199 432 201
rect 434 200 459 201
rect 434 199 444 200
rect 431 198 444 199
rect 446 198 455 200
rect 457 198 459 200
rect 431 197 459 198
rect 406 186 411 188
rect 431 187 435 197
rect 406 184 407 186
rect 409 184 411 186
rect 424 185 435 187
rect 406 182 421 184
rect 407 180 421 182
rect 424 183 425 185
rect 427 183 435 185
rect 424 181 435 183
rect 410 174 414 176
rect 410 172 411 174
rect 413 172 414 174
rect 410 166 414 172
rect 417 175 421 180
rect 455 177 459 197
rect 443 176 449 177
rect 417 174 432 175
rect 417 172 428 174
rect 430 172 432 174
rect 417 171 432 172
rect 443 174 445 176
rect 447 174 449 176
rect 443 166 449 174
rect 453 176 459 177
rect 453 174 455 176
rect 457 174 459 176
rect 453 173 459 174
rect 493 210 502 212
rect 504 210 506 212
rect 493 209 506 210
rect 481 205 497 209
rect 481 195 485 205
rect 505 201 509 203
rect 481 193 482 195
rect 484 193 485 195
rect 481 188 485 193
rect 488 192 489 198
rect 505 199 506 201
rect 508 200 533 201
rect 508 199 518 200
rect 505 198 518 199
rect 520 198 529 200
rect 531 198 533 200
rect 505 197 533 198
rect 480 186 485 188
rect 505 187 509 197
rect 480 184 481 186
rect 483 184 485 186
rect 498 185 509 187
rect 480 182 495 184
rect 481 180 495 182
rect 498 183 499 185
rect 501 183 509 185
rect 498 181 509 183
rect 484 174 488 176
rect 484 172 485 174
rect 487 172 488 174
rect 484 166 488 172
rect 491 175 495 180
rect 529 177 533 197
rect 517 176 523 177
rect 491 174 506 175
rect 491 172 502 174
rect 504 172 506 174
rect 491 171 506 172
rect 517 174 519 176
rect 521 174 523 176
rect 517 166 523 174
rect 527 176 533 177
rect 527 174 529 176
rect 531 174 533 176
rect 527 173 533 174
rect -18 149 -12 150
rect -18 147 -16 149
rect -14 147 -12 149
rect -18 146 -12 147
rect 1 149 7 150
rect 1 147 3 149
rect 5 147 7 149
rect 1 146 7 147
rect 65 144 71 150
rect 27 143 47 144
rect 27 141 43 143
rect 45 141 47 143
rect 65 142 67 144
rect 69 142 71 144
rect 65 141 71 142
rect 78 141 82 143
rect 27 140 47 141
rect -21 136 -3 137
rect -21 134 -7 136
rect -5 134 -3 136
rect -21 133 -3 134
rect -21 127 -17 133
rect -21 125 -20 127
rect -18 125 -17 127
rect -25 104 -24 115
rect -21 112 -17 125
rect -2 120 4 121
rect -21 108 -6 112
rect -10 104 -6 108
rect 15 137 16 139
rect 27 136 31 140
rect 78 139 79 141
rect 81 139 82 141
rect 19 132 31 136
rect 19 127 23 132
rect 19 125 20 127
rect 22 125 23 127
rect 19 113 23 125
rect 52 136 56 138
rect 52 134 53 136
rect 55 134 56 136
rect 52 128 56 134
rect 78 136 82 139
rect 78 132 102 136
rect 52 124 63 128
rect 19 110 36 113
rect 19 109 33 110
rect 32 108 33 109
rect 35 108 36 110
rect 21 105 27 106
rect -10 103 7 104
rect -10 101 3 103
rect 5 101 7 103
rect -10 100 7 101
rect 21 103 23 105
rect 25 103 27 105
rect -18 96 -12 97
rect -18 94 -16 96
rect -14 94 -12 96
rect 21 94 27 103
rect 32 103 36 108
rect 59 118 63 124
rect 98 128 102 132
rect 78 127 94 128
rect 78 125 90 127
rect 92 125 94 127
rect 78 124 94 125
rect 98 126 103 128
rect 98 124 100 126
rect 102 124 103 126
rect 78 118 82 124
rect 98 122 103 124
rect 98 120 102 122
rect 59 117 82 118
rect 59 115 61 117
rect 63 115 82 117
rect 59 114 82 115
rect 32 101 33 103
rect 35 101 36 103
rect 32 99 36 101
rect 41 103 47 104
rect 41 101 43 103
rect 45 101 47 103
rect 41 94 47 101
rect 70 103 74 105
rect 70 101 71 103
rect 73 101 74 103
rect 70 96 74 101
rect 78 103 82 114
rect 86 117 102 120
rect 86 115 87 117
rect 89 116 102 117
rect 89 115 90 116
rect 86 110 90 115
rect 86 108 87 110
rect 89 108 90 110
rect 86 106 90 108
rect 169 144 175 150
rect 276 149 282 150
rect 276 147 278 149
rect 280 147 282 149
rect 276 146 282 147
rect 295 149 301 150
rect 295 147 297 149
rect 299 147 301 149
rect 295 146 301 147
rect 131 143 151 144
rect 131 141 147 143
rect 149 141 151 143
rect 169 142 171 144
rect 173 142 175 144
rect 169 141 175 142
rect 182 141 186 143
rect 131 140 151 141
rect 119 137 120 139
rect 131 136 135 140
rect 182 139 183 141
rect 185 139 186 141
rect 228 143 248 144
rect 228 141 230 143
rect 232 141 248 143
rect 228 140 248 141
rect 123 132 135 136
rect 123 127 127 132
rect 123 125 124 127
rect 126 125 127 127
rect 123 113 127 125
rect 156 136 160 138
rect 156 134 157 136
rect 159 134 160 136
rect 156 128 160 134
rect 182 136 186 139
rect 182 132 206 136
rect 156 124 167 128
rect 123 110 140 113
rect 123 109 137 110
rect 136 108 137 109
rect 139 108 140 110
rect 125 105 131 106
rect 125 103 127 105
rect 129 103 131 105
rect 78 102 111 103
rect 78 100 107 102
rect 109 100 111 102
rect 78 99 111 100
rect 70 94 71 96
rect 73 94 74 96
rect 125 94 131 103
rect 136 103 140 108
rect 163 118 167 124
rect 202 128 206 132
rect 182 127 198 128
rect 182 125 194 127
rect 196 125 198 127
rect 182 124 198 125
rect 202 126 207 128
rect 202 124 204 126
rect 206 124 207 126
rect 182 118 186 124
rect 202 122 207 124
rect 202 120 206 122
rect 163 117 186 118
rect 163 115 165 117
rect 167 115 186 117
rect 163 114 186 115
rect 136 101 137 103
rect 139 101 140 103
rect 136 99 140 101
rect 145 103 151 104
rect 145 101 147 103
rect 149 101 151 103
rect 145 94 151 101
rect 174 103 178 105
rect 174 101 175 103
rect 177 101 178 103
rect 174 96 178 101
rect 182 103 186 114
rect 190 117 206 120
rect 190 115 191 117
rect 193 116 206 117
rect 193 115 194 116
rect 190 110 194 115
rect 244 136 248 140
rect 259 137 260 139
rect 244 132 256 136
rect 252 127 256 132
rect 252 125 253 127
rect 255 125 256 127
rect 190 108 191 110
rect 193 108 194 110
rect 190 106 194 108
rect 252 113 256 125
rect 336 144 340 150
rect 336 142 337 144
rect 339 142 340 144
rect 336 140 340 142
rect 343 144 358 145
rect 343 142 354 144
rect 356 142 358 144
rect 343 141 358 142
rect 369 142 375 150
rect 410 144 414 150
rect 286 136 304 137
rect 286 134 288 136
rect 290 134 304 136
rect 286 133 304 134
rect 300 127 304 133
rect 300 125 301 127
rect 303 125 304 127
rect 279 120 285 121
rect 239 110 256 113
rect 239 108 240 110
rect 242 109 256 110
rect 242 108 243 109
rect 228 103 234 104
rect 182 102 215 103
rect 182 100 211 102
rect 213 100 215 102
rect 182 99 215 100
rect 228 101 230 103
rect 232 101 234 103
rect 174 94 175 96
rect 177 94 178 96
rect 228 94 234 101
rect 239 103 243 108
rect 300 112 304 125
rect 289 108 304 112
rect 239 101 240 103
rect 242 101 243 103
rect 239 99 243 101
rect 248 105 254 106
rect 248 103 250 105
rect 252 103 254 105
rect 289 104 293 108
rect 307 104 308 115
rect 248 94 254 103
rect 276 103 293 104
rect 276 101 278 103
rect 280 101 293 103
rect 276 100 293 101
rect 343 136 347 141
rect 369 140 371 142
rect 373 140 375 142
rect 369 139 375 140
rect 379 142 385 143
rect 379 140 381 142
rect 383 140 385 142
rect 379 139 385 140
rect 333 134 347 136
rect 332 132 347 134
rect 350 133 361 135
rect 332 130 333 132
rect 335 130 337 132
rect 332 128 337 130
rect 350 131 351 133
rect 353 131 361 133
rect 350 129 361 131
rect 333 123 337 128
rect 333 121 334 123
rect 336 121 337 123
rect 333 111 337 121
rect 357 119 361 129
rect 381 119 385 139
rect 357 118 385 119
rect 357 117 370 118
rect 357 115 358 117
rect 360 116 370 117
rect 372 116 381 118
rect 383 116 385 118
rect 360 115 385 116
rect 410 142 411 144
rect 413 142 414 144
rect 410 140 414 142
rect 417 144 432 145
rect 417 142 428 144
rect 430 142 432 144
rect 417 141 432 142
rect 443 142 449 150
rect 484 144 488 150
rect 417 136 421 141
rect 443 140 445 142
rect 447 140 449 142
rect 443 139 449 140
rect 453 142 459 143
rect 453 140 455 142
rect 457 140 459 142
rect 453 139 459 140
rect 407 134 421 136
rect 406 132 421 134
rect 424 133 435 135
rect 406 130 407 132
rect 409 130 411 132
rect 406 128 411 130
rect 424 131 425 133
rect 427 131 435 133
rect 424 129 435 131
rect 357 113 361 115
rect 333 107 349 111
rect 345 106 358 107
rect 345 104 354 106
rect 356 104 358 106
rect 345 103 358 104
rect 407 123 411 128
rect 407 121 408 123
rect 410 121 411 123
rect 407 111 411 121
rect 431 119 435 129
rect 455 119 459 139
rect 431 118 459 119
rect 431 117 444 118
rect 431 115 432 117
rect 434 116 444 117
rect 446 116 455 118
rect 457 116 459 118
rect 434 115 459 116
rect 484 142 485 144
rect 487 142 488 144
rect 484 140 488 142
rect 491 144 506 145
rect 491 142 502 144
rect 504 142 506 144
rect 491 141 506 142
rect 517 142 523 150
rect 431 113 435 115
rect 407 107 423 111
rect 419 106 432 107
rect 419 104 428 106
rect 430 104 432 106
rect 419 103 432 104
rect 491 136 495 141
rect 517 140 519 142
rect 521 140 523 142
rect 517 139 523 140
rect 527 142 533 143
rect 527 140 529 142
rect 531 140 533 142
rect 527 139 533 140
rect 481 134 495 136
rect 480 132 495 134
rect 498 133 509 135
rect 480 130 481 132
rect 483 130 485 132
rect 480 128 485 130
rect 498 131 499 133
rect 501 131 509 133
rect 498 129 509 131
rect 481 123 485 128
rect 481 121 482 123
rect 484 121 485 123
rect 481 111 485 121
rect 488 118 489 124
rect 505 119 509 129
rect 529 119 533 139
rect 505 118 533 119
rect 505 117 518 118
rect 505 115 506 117
rect 508 116 518 117
rect 520 116 529 118
rect 531 116 533 118
rect 508 115 533 116
rect 505 113 509 115
rect 481 107 497 111
rect 493 106 506 107
rect 493 104 502 106
rect 504 104 506 106
rect 493 103 506 104
rect 295 96 301 97
rect 295 94 297 96
rect 299 94 301 96
rect 335 96 341 97
rect 335 94 337 96
rect 339 94 341 96
rect 370 96 374 98
rect 370 94 371 96
rect 373 94 374 96
rect 409 96 415 97
rect 409 94 411 96
rect 413 94 415 96
rect 444 96 448 98
rect 444 94 445 96
rect 447 94 448 96
rect 483 96 489 97
rect 483 94 485 96
rect 487 94 489 96
rect 518 96 522 98
rect 518 94 519 96
rect 521 94 522 96
rect -18 76 -16 78
rect -14 76 -12 78
rect -18 75 -12 76
rect -10 71 7 72
rect -10 69 3 71
rect 5 69 7 71
rect -10 68 7 69
rect 21 69 27 78
rect -25 57 -24 68
rect -10 64 -6 68
rect 21 67 23 69
rect 25 67 27 69
rect 21 66 27 67
rect 32 71 36 73
rect 32 69 33 71
rect 35 69 36 71
rect -21 60 -6 64
rect -21 47 -17 60
rect 32 64 36 69
rect 41 71 47 78
rect 70 76 71 78
rect 73 76 74 78
rect 41 69 43 71
rect 45 69 47 71
rect 41 68 47 69
rect 70 71 74 76
rect 70 69 71 71
rect 73 69 74 71
rect 70 67 74 69
rect 78 72 111 73
rect 78 70 107 72
rect 109 70 111 72
rect 78 69 111 70
rect 125 69 131 78
rect 32 63 33 64
rect 19 62 33 63
rect 35 62 36 64
rect 19 59 36 62
rect -2 51 4 52
rect -21 45 -20 47
rect -18 45 -17 47
rect -21 39 -17 45
rect -21 38 -3 39
rect -21 36 -7 38
rect -5 36 -3 38
rect -21 35 -3 36
rect 19 47 23 59
rect 78 58 82 69
rect 125 67 127 69
rect 129 67 131 69
rect 125 66 131 67
rect 136 71 140 73
rect 136 69 137 71
rect 139 69 140 71
rect 59 57 82 58
rect 59 55 61 57
rect 63 55 82 57
rect 59 54 82 55
rect 59 48 63 54
rect 19 45 20 47
rect 22 45 23 47
rect 19 40 23 45
rect 19 36 31 40
rect 15 33 16 35
rect 27 32 31 36
rect 52 44 63 48
rect 52 38 56 44
rect 78 48 82 54
rect 86 64 90 66
rect 86 62 87 64
rect 89 62 90 64
rect 86 57 90 62
rect 86 55 87 57
rect 89 56 90 57
rect 89 55 102 56
rect 86 52 102 55
rect 98 50 102 52
rect 98 48 103 50
rect 78 47 94 48
rect 78 45 90 47
rect 92 45 94 47
rect 78 44 94 45
rect 98 46 100 48
rect 102 46 103 48
rect 98 44 103 46
rect 52 36 53 38
rect 55 36 56 38
rect 52 34 56 36
rect 98 40 102 44
rect 78 36 102 40
rect 78 33 82 36
rect 27 31 47 32
rect 78 31 79 33
rect 81 31 82 33
rect 27 29 43 31
rect 45 29 47 31
rect 27 28 47 29
rect 65 30 71 31
rect 65 28 67 30
rect 69 28 71 30
rect 78 29 82 31
rect 136 64 140 69
rect 145 71 151 78
rect 174 76 175 78
rect 177 76 178 78
rect 145 69 147 71
rect 149 69 151 71
rect 145 68 151 69
rect 174 71 178 76
rect 174 69 175 71
rect 177 69 178 71
rect 174 67 178 69
rect 182 72 215 73
rect 182 70 211 72
rect 213 70 215 72
rect 182 69 215 70
rect 228 71 234 78
rect 228 69 230 71
rect 232 69 234 71
rect 136 63 137 64
rect 123 62 137 63
rect 139 62 140 64
rect 123 59 140 62
rect 123 47 127 59
rect 182 58 186 69
rect 228 68 234 69
rect 239 71 243 73
rect 239 69 240 71
rect 242 69 243 71
rect 163 57 186 58
rect 163 55 165 57
rect 167 55 186 57
rect 163 54 186 55
rect 163 48 167 54
rect 123 45 124 47
rect 126 45 127 47
rect 123 40 127 45
rect 123 36 135 40
rect 119 33 120 35
rect -18 25 -12 26
rect -18 23 -16 25
rect -14 23 -12 25
rect -18 22 -12 23
rect 1 25 7 26
rect 1 23 3 25
rect 5 23 7 25
rect 1 22 7 23
rect 65 22 71 28
rect 131 32 135 36
rect 156 44 167 48
rect 156 38 160 44
rect 182 48 186 54
rect 190 64 194 66
rect 190 62 191 64
rect 193 62 194 64
rect 190 57 194 62
rect 190 55 191 57
rect 193 56 194 57
rect 193 55 206 56
rect 190 52 206 55
rect 202 50 206 52
rect 202 48 207 50
rect 182 47 198 48
rect 182 45 194 47
rect 196 45 198 47
rect 182 44 198 45
rect 202 46 204 48
rect 206 46 207 48
rect 202 44 207 46
rect 156 36 157 38
rect 159 36 160 38
rect 156 34 160 36
rect 202 40 206 44
rect 182 36 206 40
rect 239 64 243 69
rect 248 69 254 78
rect 295 76 297 78
rect 299 76 301 78
rect 295 75 301 76
rect 335 76 337 78
rect 339 76 341 78
rect 335 75 341 76
rect 370 76 371 78
rect 373 76 374 78
rect 370 74 374 76
rect 409 76 411 78
rect 413 76 415 78
rect 409 75 415 76
rect 444 76 445 78
rect 447 76 448 78
rect 444 74 448 76
rect 483 76 485 78
rect 487 76 489 78
rect 483 75 489 76
rect 518 76 519 78
rect 521 76 522 78
rect 518 74 522 76
rect 248 67 250 69
rect 252 67 254 69
rect 276 71 293 72
rect 276 69 278 71
rect 280 69 293 71
rect 276 68 293 69
rect 248 66 254 67
rect 239 62 240 64
rect 242 63 243 64
rect 242 62 256 63
rect 239 59 256 62
rect 182 33 186 36
rect 131 31 151 32
rect 182 31 183 33
rect 185 31 186 33
rect 252 47 256 59
rect 252 45 253 47
rect 255 45 256 47
rect 252 40 256 45
rect 244 36 256 40
rect 289 64 293 68
rect 289 60 304 64
rect 279 51 285 52
rect 244 32 248 36
rect 259 33 260 35
rect 300 47 304 60
rect 307 57 308 68
rect 300 45 301 47
rect 303 45 304 47
rect 300 39 304 45
rect 286 38 304 39
rect 286 36 288 38
rect 290 36 304 38
rect 286 35 304 36
rect 345 68 358 69
rect 345 66 354 68
rect 356 66 358 68
rect 345 65 358 66
rect 333 61 349 65
rect 333 51 337 61
rect 419 68 432 69
rect 357 57 361 59
rect 333 49 334 51
rect 336 49 337 51
rect 333 44 337 49
rect 332 42 337 44
rect 357 55 358 57
rect 360 56 385 57
rect 360 55 370 56
rect 357 54 370 55
rect 372 54 381 56
rect 383 54 385 56
rect 357 53 385 54
rect 357 43 361 53
rect 332 40 333 42
rect 335 40 337 42
rect 350 41 361 43
rect 332 38 347 40
rect 333 36 347 38
rect 350 39 351 41
rect 353 39 361 41
rect 350 37 361 39
rect 131 29 147 31
rect 149 29 151 31
rect 131 28 151 29
rect 169 30 175 31
rect 169 28 171 30
rect 173 28 175 30
rect 182 29 186 31
rect 228 31 248 32
rect 228 29 230 31
rect 232 29 248 31
rect 228 28 248 29
rect 169 22 175 28
rect 336 30 340 32
rect 336 28 337 30
rect 339 28 340 30
rect 276 25 282 26
rect 276 23 278 25
rect 280 23 282 25
rect 276 22 282 23
rect 295 25 301 26
rect 295 23 297 25
rect 299 23 301 25
rect 295 22 301 23
rect 336 22 340 28
rect 343 31 347 36
rect 381 33 385 53
rect 369 32 375 33
rect 343 30 358 31
rect 343 28 354 30
rect 356 28 358 30
rect 343 27 358 28
rect 369 30 371 32
rect 373 30 375 32
rect 369 22 375 30
rect 379 32 385 33
rect 379 30 381 32
rect 383 30 385 32
rect 379 29 385 30
rect 419 66 428 68
rect 430 66 432 68
rect 419 65 432 66
rect 407 61 423 65
rect 407 51 411 61
rect 493 68 506 69
rect 431 57 435 59
rect 407 49 408 51
rect 410 49 411 51
rect 407 44 411 49
rect 431 55 432 57
rect 434 56 459 57
rect 434 55 444 56
rect 431 54 444 55
rect 446 54 455 56
rect 457 54 459 56
rect 431 53 459 54
rect 406 42 411 44
rect 431 43 435 53
rect 406 40 407 42
rect 409 40 411 42
rect 424 41 435 43
rect 406 38 421 40
rect 407 36 421 38
rect 424 39 425 41
rect 427 39 435 41
rect 424 37 435 39
rect 410 30 414 32
rect 410 28 411 30
rect 413 28 414 30
rect 410 22 414 28
rect 417 31 421 36
rect 455 33 459 53
rect 443 32 449 33
rect 417 30 432 31
rect 417 28 428 30
rect 430 28 432 30
rect 417 27 432 28
rect 443 30 445 32
rect 447 30 449 32
rect 443 22 449 30
rect 453 32 459 33
rect 453 30 455 32
rect 457 30 459 32
rect 453 29 459 30
rect 493 66 502 68
rect 504 66 506 68
rect 493 65 506 66
rect 481 61 497 65
rect 481 51 485 61
rect 505 57 509 59
rect 481 49 482 51
rect 484 49 485 51
rect 481 44 485 49
rect 488 48 489 54
rect 505 55 506 57
rect 508 56 533 57
rect 508 55 518 56
rect 505 54 518 55
rect 520 54 529 56
rect 531 54 533 56
rect 505 53 533 54
rect 480 42 485 44
rect 505 43 509 53
rect 480 40 481 42
rect 483 40 485 42
rect 498 41 509 43
rect 480 38 495 40
rect 481 36 495 38
rect 498 39 499 41
rect 501 39 509 41
rect 498 37 509 39
rect 484 30 488 32
rect 484 28 485 30
rect 487 28 488 30
rect 484 22 488 28
rect 491 31 495 36
rect 529 33 533 53
rect 517 32 523 33
rect 491 30 506 31
rect 491 28 502 30
rect 504 28 506 30
rect 491 27 506 28
rect 517 30 519 32
rect 521 30 523 32
rect 517 22 523 30
rect 527 32 533 33
rect 527 30 529 32
rect 531 30 533 32
rect 527 29 533 30
<< via1 >>
rect 4 269 6 271
rect 4 256 6 258
rect 36 278 38 280
rect 12 256 14 258
rect 61 278 63 280
rect 69 278 71 280
rect 44 254 46 256
rect 53 254 55 256
rect 108 261 110 263
rect 116 269 118 271
rect 140 278 142 280
rect 131 269 133 271
rect 165 278 167 280
rect 139 261 141 263
rect 148 254 150 256
rect 212 273 214 275
rect 157 254 159 256
rect 237 278 239 280
rect 229 261 231 263
rect 277 278 279 280
rect 261 264 263 266
rect 277 261 279 263
rect 309 263 311 265
rect 326 271 328 273
rect 341 261 343 263
rect 368 271 370 273
rect 400 267 402 269
rect 417 269 419 271
rect 490 267 492 269
rect 516 276 518 278
rect -28 214 -26 216
rect 4 202 6 204
rect 12 202 14 204
rect 44 204 46 206
rect 4 189 6 191
rect 53 204 55 206
rect 36 180 38 182
rect 108 197 110 199
rect 61 180 63 182
rect 148 204 150 206
rect 116 189 118 191
rect 139 197 141 199
rect 157 204 159 206
rect 131 189 133 191
rect 140 180 142 182
rect 165 180 167 182
rect 229 197 231 199
rect 212 185 214 187
rect 236 180 238 182
rect 277 197 279 199
rect 261 194 263 196
rect 309 195 311 197
rect 277 180 279 182
rect 326 187 328 189
rect 341 197 343 199
rect 368 187 370 189
rect 400 191 402 193
rect 417 189 419 191
rect 490 191 492 193
rect 516 182 518 184
rect -36 131 -34 133
rect 4 125 6 127
rect 4 112 6 114
rect 36 134 38 136
rect 12 112 14 114
rect 61 134 63 136
rect 69 134 71 136
rect 44 117 46 119
rect 44 109 46 111
rect 52 109 54 111
rect 108 117 110 119
rect 116 125 118 127
rect 140 134 142 136
rect 131 125 133 127
rect 165 134 167 136
rect 139 117 141 119
rect 148 110 150 112
rect 212 129 214 131
rect 157 110 159 112
rect 237 134 239 136
rect 229 117 231 119
rect 277 134 279 136
rect 261 120 263 122
rect 277 117 279 119
rect 309 119 311 121
rect 326 127 328 129
rect 341 117 343 119
rect 368 127 370 129
rect 400 123 402 125
rect 417 125 419 127
rect 490 123 492 125
rect 516 132 518 134
rect -28 47 -26 49
rect 4 58 6 60
rect 12 58 14 60
rect 44 60 46 62
rect 4 45 6 47
rect 53 60 55 62
rect 36 36 38 38
rect 108 53 110 55
rect 61 36 63 38
rect 148 60 150 62
rect 116 45 118 47
rect 139 53 141 55
rect 157 60 159 62
rect 140 36 142 38
rect 165 36 167 38
rect 229 61 231 63
rect 212 41 214 43
rect 237 45 239 47
rect 277 61 279 63
rect 261 50 263 52
rect 277 45 279 47
rect 309 51 311 53
rect 326 43 328 45
rect 341 53 343 55
rect 368 43 370 45
rect 400 47 402 49
rect 417 45 419 47
rect 490 47 492 49
rect 516 38 518 40
<< via2 >>
rect 69 278 71 280
rect 237 278 239 280
rect 277 278 279 280
rect 131 269 133 271
rect 53 254 55 256
rect 229 261 231 263
rect 277 261 279 263
rect -28 214 -26 216
rect 53 204 55 206
rect 131 189 133 191
rect 229 197 231 199
rect 277 197 279 199
rect 61 180 63 182
rect 236 180 238 182
rect 277 180 279 182
rect -36 145 -34 147
rect 69 134 71 136
rect 237 134 239 136
rect 277 134 279 136
rect 131 125 133 127
rect 44 117 46 119
rect 229 117 231 119
rect 277 117 279 119
rect 44 60 46 62
rect -28 47 -26 49
rect 229 61 231 63
rect 277 61 279 63
rect 237 45 239 47
rect 277 45 279 47
<< labels >>
rlabel polyct1 382 66 382 66 1 s0
rlabel polyct1 456 66 456 66 1 s0
rlabel polyct1 530 66 530 66 1 s1
rlabel alu1 383 83 383 83 1 vdd!
rlabel alu1 501 17 501 17 1 vss!
rlabel pwell 211 40 215 44 1 sum0
rlabel alu1 473 48 477 51 1 aluout0
rlabel polyct1 382 106 382 106 5 s0
rlabel polyct1 456 106 456 106 5 s0
rlabel polyct1 530 106 530 106 5 s1
rlabel alu1 383 89 383 89 5 vdd!
rlabel alu1 501 155 501 155 5 vss!
rlabel pwell 211 128 215 132 1 sum1
rlabel alu1 473 119 477 122 1 aluout1
rlabel polyct1 382 210 382 210 1 s0
rlabel polyct1 456 210 456 210 1 s0
rlabel polyct1 530 210 530 210 1 s1
rlabel alu1 383 227 383 227 1 vdd!
rlabel alu1 501 161 501 161 1 vss!
rlabel polyct1 382 250 382 250 5 s0
rlabel polyct1 456 250 456 250 5 s0
rlabel polyct1 530 250 530 250 5 s1
rlabel alu1 383 233 383 233 5 vdd!
rlabel alu1 501 299 501 299 5 vss!
rlabel pwell 211 184 215 188 1 sum2
rlabel alu1 473 192 477 196 1 aluout2
rlabel alu1 473 263 477 266 1 aluout3
rlabel pwell 211 272 215 276 1 sum3
rlabel alu1 36 130 38 130 1 a1
rlabel alu1 -27 274 -27 274 1 cout
rlabel alu1 37 274 37 274 1 a3
rlabel alu1 140 43 140 43 1 cin0
rlabel alu2 48 181 48 181 1 a2
rlabel alu2 49 255 49 255 1 b3
rlabel alu2 49 205 49 205 1 b2
rlabel alu2 49 110 49 110 1 b1
rlabel alu3 49 61 49 61 1 b0
rlabel alu1 140 129 140 129 1 cin1
rlabel alu3 -28 144 -28 144 3 cout1
rlabel alu1 -28 44 -28 44 1 cout0
rlabel alu2 25 46 25 46 1 a0
rlabel alu3 240 46 240 46 1 a0
<< end >>
