magic
tech scmos
timestamp 1636182940
<< ab >>
rect 2 55 52 104
rect 2 52 40 55
rect 44 52 52 55
rect 2 4 52 52
rect 76 55 126 104
rect 76 53 115 55
rect 117 53 126 55
rect 76 4 126 53
rect 153 84 397 92
rect 153 68 233 84
rect 153 67 228 68
rect 230 67 233 68
rect 153 52 233 67
rect 234 52 337 84
rect 338 52 401 84
rect 153 51 212 52
rect 214 51 401 52
rect 153 48 401 51
rect 153 47 252 48
rect 253 47 401 48
rect 153 28 401 47
rect 156 20 399 28
rect 228 15 234 20
rect 332 15 338 20
rect 423 4 573 104
<< nwell >>
rect 0 52 575 108
<< pwell >>
rect 0 0 575 52
<< poly >>
rect 37 99 39 103
rect 111 99 113 103
rect 448 99 450 103
rect 460 99 462 103
rect 472 99 474 103
rect 480 99 482 103
rect 492 99 494 103
rect 504 99 506 103
rect 512 99 514 103
rect 536 99 538 103
rect 548 99 550 103
rect 13 89 15 93
rect 25 89 27 93
rect 13 67 15 69
rect 9 65 15 67
rect 9 63 11 65
rect 13 63 15 65
rect 9 61 15 63
rect 25 57 27 69
rect 91 89 93 93
rect 99 89 101 93
rect 175 86 177 90
rect 182 86 184 90
rect 162 76 164 81
rect 25 55 33 57
rect 25 53 29 55
rect 31 53 33 55
rect 25 51 33 53
rect 9 45 15 47
rect 9 43 11 45
rect 13 43 15 45
rect 9 41 15 43
rect 19 45 25 47
rect 37 45 39 59
rect 91 57 93 59
rect 87 55 93 57
rect 99 57 101 59
rect 99 55 107 57
rect 87 47 89 55
rect 99 53 103 55
rect 105 53 107 55
rect 99 51 107 53
rect 19 43 21 45
rect 23 43 39 45
rect 19 41 25 43
rect 13 39 15 41
rect 25 35 33 37
rect 25 33 29 35
rect 31 33 33 35
rect 25 31 33 33
rect 25 29 27 31
rect 37 29 39 43
rect 83 45 89 47
rect 83 43 85 45
rect 87 43 89 45
rect 83 41 89 43
rect 93 45 99 47
rect 111 45 113 59
rect 250 86 252 90
rect 202 77 204 81
rect 212 79 214 84
rect 222 79 224 84
rect 162 55 164 58
rect 175 55 177 65
rect 182 62 184 65
rect 182 60 188 62
rect 182 58 184 60
rect 186 58 188 60
rect 182 56 188 58
rect 162 53 168 55
rect 162 51 164 53
rect 166 51 168 53
rect 162 49 168 51
rect 172 53 178 55
rect 172 51 174 53
rect 176 51 178 53
rect 172 49 178 51
rect 162 46 164 49
rect 172 46 174 49
rect 182 46 184 56
rect 202 55 204 59
rect 212 55 214 66
rect 222 63 224 66
rect 222 61 228 63
rect 222 59 224 61
rect 226 59 228 61
rect 222 57 228 59
rect 235 61 241 63
rect 235 59 237 61
rect 239 59 241 61
rect 286 86 288 90
rect 266 77 268 81
rect 276 77 278 81
rect 354 86 356 90
rect 306 77 308 81
rect 316 79 318 84
rect 326 79 328 84
rect 235 57 241 59
rect 202 53 208 55
rect 202 51 204 53
rect 206 51 208 53
rect 202 49 208 51
rect 212 53 218 55
rect 212 51 214 53
rect 216 51 218 53
rect 212 49 218 51
rect 93 43 95 45
rect 97 43 113 45
rect 93 41 99 43
rect 87 29 89 41
rect 99 35 107 37
rect 99 33 103 35
rect 105 33 107 35
rect 99 31 107 33
rect 99 29 101 31
rect 111 29 113 43
rect 202 44 204 49
rect 215 44 217 49
rect 222 44 224 57
rect 239 56 241 57
rect 250 56 252 59
rect 266 56 268 59
rect 239 54 252 56
rect 258 54 268 56
rect 276 55 278 59
rect 286 56 288 59
rect 242 46 244 54
rect 258 50 260 54
rect 251 48 260 50
rect 272 53 278 55
rect 272 51 274 53
rect 276 51 278 53
rect 272 49 278 51
rect 282 54 288 56
rect 282 52 284 54
rect 286 52 288 54
rect 282 50 288 52
rect 306 55 308 59
rect 316 55 318 66
rect 326 63 328 66
rect 326 61 332 63
rect 326 59 328 61
rect 330 59 332 61
rect 326 57 332 59
rect 339 61 345 63
rect 339 59 341 61
rect 343 59 345 61
rect 390 86 392 90
rect 370 77 372 81
rect 380 77 382 81
rect 436 73 438 77
rect 339 57 345 59
rect 306 53 312 55
rect 306 51 308 53
rect 310 51 312 53
rect 251 46 253 48
rect 255 46 260 48
rect 162 32 164 37
rect 172 35 174 40
rect 182 35 184 40
rect 13 15 15 19
rect 87 15 89 19
rect 99 15 101 19
rect 202 31 204 35
rect 251 44 260 46
rect 276 46 278 49
rect 258 41 260 44
rect 268 41 270 45
rect 276 44 280 46
rect 278 41 280 44
rect 285 41 287 50
rect 306 49 312 51
rect 316 53 322 55
rect 316 51 318 53
rect 320 51 322 53
rect 316 49 322 51
rect 306 44 308 49
rect 319 44 321 49
rect 326 44 328 57
rect 343 56 345 57
rect 354 56 356 59
rect 370 56 372 59
rect 343 54 356 56
rect 362 54 372 56
rect 380 55 382 59
rect 390 56 392 59
rect 436 57 438 59
rect 346 46 348 54
rect 362 50 364 54
rect 355 48 364 50
rect 376 53 382 55
rect 376 51 378 53
rect 380 51 382 53
rect 376 49 382 51
rect 386 54 392 56
rect 386 52 388 54
rect 390 52 392 54
rect 386 50 392 52
rect 428 55 438 57
rect 428 53 430 55
rect 432 53 438 55
rect 428 51 438 53
rect 355 46 357 48
rect 359 46 364 48
rect 242 34 244 37
rect 215 28 217 33
rect 222 28 224 33
rect 242 32 247 34
rect 245 24 247 32
rect 258 28 260 32
rect 268 24 270 32
rect 306 31 308 35
rect 355 44 364 46
rect 380 46 382 49
rect 362 41 364 44
rect 372 41 374 45
rect 380 44 384 46
rect 382 41 384 44
rect 389 41 391 50
rect 436 41 438 51
rect 448 57 450 79
rect 460 77 462 79
rect 454 75 462 77
rect 454 73 456 75
rect 458 73 462 75
rect 454 71 462 73
rect 448 55 456 57
rect 448 53 452 55
rect 454 53 456 55
rect 448 51 456 53
rect 346 34 348 37
rect 278 24 280 29
rect 285 24 287 29
rect 245 22 270 24
rect 319 28 321 33
rect 326 28 328 33
rect 346 32 351 34
rect 349 24 351 32
rect 362 28 364 32
rect 372 24 374 32
rect 382 24 384 29
rect 389 24 391 29
rect 349 22 374 24
rect 436 29 438 33
rect 448 27 450 51
rect 460 45 462 71
rect 472 67 474 79
rect 468 65 474 67
rect 468 63 470 65
rect 472 63 474 65
rect 468 61 474 63
rect 470 55 476 57
rect 480 55 482 79
rect 492 77 494 79
rect 504 77 506 79
rect 470 53 472 55
rect 474 53 482 55
rect 470 51 476 53
rect 460 43 474 45
rect 454 35 462 37
rect 454 33 456 35
rect 458 33 462 35
rect 454 31 462 33
rect 460 27 462 31
rect 472 27 474 43
rect 480 27 482 53
rect 490 75 494 77
rect 500 75 506 77
rect 490 37 492 75
rect 500 57 502 75
rect 512 67 514 79
rect 524 73 526 76
rect 506 65 514 67
rect 506 63 508 65
rect 510 63 514 65
rect 506 61 514 63
rect 560 79 562 83
rect 496 55 502 57
rect 524 55 526 59
rect 496 53 498 55
rect 500 53 526 55
rect 496 51 502 53
rect 500 43 502 51
rect 486 35 492 37
rect 486 33 488 35
rect 490 33 492 35
rect 486 31 492 33
rect 496 41 502 43
rect 506 45 514 47
rect 506 43 508 45
rect 510 43 514 45
rect 506 41 514 43
rect 524 41 526 53
rect 536 47 538 59
rect 548 47 550 59
rect 560 57 562 59
rect 554 55 562 57
rect 554 53 556 55
rect 558 53 560 55
rect 554 51 560 53
rect 564 47 570 49
rect 536 45 566 47
rect 568 45 570 47
rect 496 27 498 41
rect 502 35 508 37
rect 502 33 504 35
rect 506 33 508 35
rect 502 31 508 33
rect 492 25 498 27
rect 492 23 494 25
rect 504 23 506 31
rect 512 23 514 41
rect 524 30 526 33
rect 536 31 538 45
rect 548 31 550 45
rect 564 43 570 45
rect 554 37 560 39
rect 554 35 556 37
rect 558 35 560 37
rect 554 33 562 35
rect 560 31 562 33
rect 448 11 450 15
rect 460 11 462 15
rect 472 11 474 15
rect 480 11 482 15
rect 560 17 562 21
rect 25 5 27 9
rect 37 5 39 9
rect 111 5 113 9
rect 492 7 494 11
rect 504 7 506 11
rect 512 7 514 11
rect 536 7 538 11
rect 548 7 550 11
<< ndif >>
rect 5 25 13 39
rect 5 23 7 25
rect 9 23 13 25
rect 5 19 13 23
rect 15 29 23 39
rect 155 44 162 46
rect 155 42 157 44
rect 159 42 162 44
rect 155 40 162 42
rect 157 37 162 40
rect 164 40 172 46
rect 174 44 182 46
rect 174 42 177 44
rect 179 42 182 44
rect 174 40 182 42
rect 184 40 191 46
rect 235 44 242 46
rect 197 41 202 44
rect 164 37 170 40
rect 166 33 170 37
rect 186 33 191 40
rect 195 39 202 41
rect 195 37 197 39
rect 199 37 202 39
rect 195 35 202 37
rect 204 35 215 44
rect 166 31 172 33
rect 166 29 168 31
rect 170 29 172 31
rect 15 19 25 29
rect 17 9 25 19
rect 27 15 37 29
rect 27 13 31 15
rect 33 13 37 15
rect 27 9 37 13
rect 39 25 47 29
rect 39 23 43 25
rect 45 23 47 25
rect 39 9 47 23
rect 79 19 87 29
rect 89 25 99 29
rect 89 23 93 25
rect 95 23 99 25
rect 89 19 99 23
rect 101 19 111 29
rect 79 15 85 19
rect 103 15 111 19
rect 79 13 81 15
rect 83 13 85 15
rect 79 11 85 13
rect 103 13 105 15
rect 107 13 111 15
rect 103 9 111 13
rect 113 25 121 29
rect 113 23 117 25
rect 119 23 121 25
rect 166 27 172 29
rect 185 31 191 33
rect 206 33 215 35
rect 217 33 222 44
rect 224 39 229 44
rect 235 42 237 44
rect 239 42 242 44
rect 235 40 242 42
rect 224 37 231 39
rect 237 37 242 40
rect 244 41 249 46
rect 339 44 346 46
rect 301 41 306 44
rect 244 37 258 41
rect 224 35 227 37
rect 229 35 231 37
rect 224 33 231 35
rect 249 36 258 37
rect 249 34 251 36
rect 253 34 258 36
rect 185 29 187 31
rect 189 29 191 31
rect 185 27 191 29
rect 206 27 213 33
rect 249 32 258 34
rect 260 39 268 41
rect 260 37 263 39
rect 265 37 268 39
rect 260 32 268 37
rect 270 37 278 41
rect 270 35 273 37
rect 275 35 278 37
rect 270 32 278 35
rect 206 25 208 27
rect 210 25 213 27
rect 206 23 213 25
rect 273 29 278 32
rect 280 29 285 41
rect 287 29 295 41
rect 299 39 306 41
rect 299 37 301 39
rect 303 37 306 39
rect 299 35 306 37
rect 308 35 319 44
rect 310 33 319 35
rect 321 33 326 44
rect 328 39 333 44
rect 339 42 341 44
rect 343 42 346 44
rect 339 40 346 42
rect 328 37 335 39
rect 341 37 346 40
rect 348 41 353 46
rect 348 37 362 41
rect 328 35 331 37
rect 333 35 335 37
rect 328 33 335 35
rect 353 36 362 37
rect 353 34 355 36
rect 357 34 362 36
rect 289 27 295 29
rect 289 25 291 27
rect 293 25 295 27
rect 113 9 121 23
rect 289 23 295 25
rect 310 27 317 33
rect 353 32 362 34
rect 364 39 372 41
rect 364 37 367 39
rect 369 37 372 39
rect 364 32 372 37
rect 374 37 382 41
rect 374 35 377 37
rect 379 35 382 37
rect 374 32 382 35
rect 310 25 312 27
rect 314 25 317 27
rect 310 23 317 25
rect 377 29 382 32
rect 384 29 389 41
rect 391 29 399 41
rect 393 27 399 29
rect 393 25 395 27
rect 397 25 399 27
rect 393 23 399 25
rect 428 33 436 41
rect 438 37 446 41
rect 438 35 442 37
rect 444 35 446 37
rect 438 33 446 35
rect 428 25 434 33
rect 464 35 470 37
rect 464 33 466 35
rect 468 33 470 35
rect 464 27 470 33
rect 428 23 430 25
rect 432 23 434 25
rect 428 21 434 23
rect 440 25 448 27
rect 440 23 442 25
rect 444 23 448 25
rect 440 15 448 23
rect 450 15 460 27
rect 462 15 472 27
rect 474 15 480 27
rect 482 25 490 27
rect 482 23 486 25
rect 488 23 490 25
rect 516 39 524 41
rect 516 37 518 39
rect 520 37 524 39
rect 516 33 524 37
rect 526 33 534 41
rect 528 31 534 33
rect 540 35 546 37
rect 540 33 542 35
rect 544 33 546 35
rect 540 31 546 33
rect 516 25 522 27
rect 516 23 518 25
rect 520 23 522 25
rect 482 15 492 23
rect 484 11 492 15
rect 494 15 504 23
rect 494 13 498 15
rect 500 13 504 15
rect 494 11 504 13
rect 506 11 512 23
rect 514 11 522 23
rect 528 15 536 31
rect 528 13 530 15
rect 532 13 536 15
rect 528 11 536 13
rect 538 11 548 31
rect 550 21 560 31
rect 562 27 570 31
rect 562 25 566 27
rect 568 25 570 27
rect 562 21 570 25
rect 550 15 558 21
rect 550 13 554 15
rect 556 13 558 15
rect 550 11 558 13
<< pdif >>
rect 5 95 11 97
rect 5 93 7 95
rect 9 93 11 95
rect 29 95 37 99
rect 29 93 31 95
rect 33 93 37 95
rect 5 89 11 93
rect 29 89 37 93
rect 5 85 13 89
rect 5 83 7 85
rect 9 83 13 85
rect 5 69 13 83
rect 15 85 25 89
rect 15 83 19 85
rect 21 83 25 85
rect 15 69 25 83
rect 27 69 37 89
rect 29 59 37 69
rect 39 85 47 99
rect 103 95 111 99
rect 103 93 105 95
rect 107 93 111 95
rect 103 89 111 93
rect 39 83 43 85
rect 45 83 47 85
rect 39 75 47 83
rect 39 73 43 75
rect 45 73 47 75
rect 39 65 47 73
rect 39 63 43 65
rect 45 63 47 65
rect 39 59 47 63
rect 79 85 91 89
rect 79 83 81 85
rect 83 83 91 85
rect 79 59 91 83
rect 93 59 99 89
rect 101 59 111 89
rect 113 85 121 99
rect 113 83 117 85
rect 119 83 121 85
rect 166 84 175 86
rect 113 75 121 83
rect 166 82 168 84
rect 170 82 175 84
rect 166 76 175 82
rect 113 73 117 75
rect 119 73 121 75
rect 113 65 121 73
rect 113 63 117 65
rect 119 63 121 65
rect 155 74 162 76
rect 155 72 157 74
rect 159 72 162 74
rect 155 67 162 72
rect 155 65 157 67
rect 159 65 162 67
rect 155 63 162 65
rect 113 59 121 63
rect 157 58 162 63
rect 164 65 175 76
rect 177 65 182 86
rect 184 79 189 86
rect 184 77 191 79
rect 206 77 212 79
rect 184 75 187 77
rect 189 75 191 77
rect 184 73 191 75
rect 184 65 189 73
rect 197 72 202 77
rect 195 70 202 72
rect 195 68 197 70
rect 199 68 202 70
rect 164 58 172 65
rect 195 63 202 68
rect 195 61 197 63
rect 199 61 202 63
rect 195 59 202 61
rect 204 75 212 77
rect 204 73 207 75
rect 209 73 212 75
rect 204 66 212 73
rect 214 77 222 79
rect 214 75 217 77
rect 219 75 222 77
rect 214 70 222 75
rect 214 68 217 70
rect 219 68 222 70
rect 214 66 222 68
rect 224 77 231 79
rect 224 75 227 77
rect 229 75 231 77
rect 224 66 231 75
rect 204 59 210 66
rect 245 65 250 86
rect 243 63 250 65
rect 243 61 245 63
rect 247 61 250 63
rect 243 59 250 61
rect 252 84 264 86
rect 252 82 255 84
rect 257 82 264 84
rect 252 77 264 82
rect 281 77 286 86
rect 252 75 255 77
rect 257 75 266 77
rect 252 59 266 75
rect 268 70 276 77
rect 268 68 271 70
rect 273 68 276 70
rect 268 63 276 68
rect 268 61 271 63
rect 273 61 276 63
rect 268 59 276 61
rect 278 70 286 77
rect 278 68 281 70
rect 283 68 286 70
rect 278 59 286 68
rect 288 80 293 86
rect 288 78 295 80
rect 288 76 291 78
rect 293 76 295 78
rect 310 77 316 79
rect 288 74 295 76
rect 288 59 293 74
rect 301 72 306 77
rect 299 70 306 72
rect 299 68 301 70
rect 303 68 306 70
rect 299 63 306 68
rect 299 61 301 63
rect 303 61 306 63
rect 299 59 306 61
rect 308 75 316 77
rect 308 73 311 75
rect 313 73 316 75
rect 308 66 316 73
rect 318 77 326 79
rect 318 75 321 77
rect 323 75 326 77
rect 318 70 326 75
rect 318 68 321 70
rect 323 68 326 70
rect 318 66 326 68
rect 328 77 335 79
rect 328 75 331 77
rect 333 75 335 77
rect 328 66 335 75
rect 308 59 314 66
rect 349 65 354 86
rect 347 63 354 65
rect 347 61 349 63
rect 351 61 354 63
rect 347 59 354 61
rect 356 84 368 86
rect 356 82 359 84
rect 361 82 368 84
rect 356 77 368 82
rect 385 77 390 86
rect 356 75 359 77
rect 361 75 370 77
rect 356 59 370 75
rect 372 70 380 77
rect 372 68 375 70
rect 377 68 380 70
rect 372 63 380 68
rect 372 61 375 63
rect 377 61 380 63
rect 372 59 380 61
rect 382 70 390 77
rect 382 68 385 70
rect 387 68 390 70
rect 382 59 390 68
rect 392 80 397 86
rect 428 85 434 87
rect 428 83 430 85
rect 432 83 434 85
rect 392 78 399 80
rect 392 76 395 78
rect 397 76 399 78
rect 392 74 399 76
rect 392 59 397 74
rect 428 73 434 83
rect 440 85 448 99
rect 440 83 442 85
rect 444 83 448 85
rect 440 79 448 83
rect 450 79 460 99
rect 462 79 472 99
rect 474 79 480 99
rect 482 85 492 99
rect 482 83 486 85
rect 488 83 492 85
rect 482 79 492 83
rect 494 95 504 99
rect 494 93 498 95
rect 500 93 504 95
rect 494 79 504 93
rect 506 79 512 99
rect 514 85 522 99
rect 514 83 518 85
rect 520 83 522 85
rect 514 79 522 83
rect 528 97 536 99
rect 528 95 530 97
rect 532 95 536 97
rect 428 59 436 73
rect 438 65 446 73
rect 438 63 442 65
rect 444 63 446 65
rect 438 59 446 63
rect 464 75 470 79
rect 464 73 466 75
rect 468 73 470 75
rect 464 71 470 73
rect 528 73 536 95
rect 516 65 524 73
rect 516 63 518 65
rect 520 63 524 65
rect 516 59 524 63
rect 526 59 536 73
rect 538 85 548 99
rect 538 83 542 85
rect 544 83 548 85
rect 538 75 548 83
rect 538 73 542 75
rect 544 73 548 75
rect 538 65 548 73
rect 538 63 542 65
rect 544 63 548 65
rect 538 59 548 63
rect 550 97 558 99
rect 550 95 554 97
rect 556 95 558 97
rect 550 85 558 95
rect 550 83 554 85
rect 556 83 558 85
rect 550 79 558 83
rect 550 75 560 79
rect 550 73 554 75
rect 556 73 560 75
rect 550 65 560 73
rect 550 63 554 65
rect 556 63 560 65
rect 550 59 560 63
rect 562 75 570 79
rect 562 73 566 75
rect 568 73 570 75
rect 562 65 570 73
rect 562 63 566 65
rect 568 63 570 65
rect 562 59 570 63
<< alu1 >>
rect 0 99 575 104
rect 0 97 81 99
rect 83 97 93 99
rect 95 97 566 99
rect 568 97 575 99
rect 0 95 530 97
rect 532 95 554 97
rect 556 95 575 97
rect 0 93 7 95
rect 9 93 31 95
rect 33 93 105 95
rect 107 93 498 95
rect 500 93 575 95
rect 0 92 575 93
rect 6 85 10 92
rect 156 87 397 92
rect 6 83 7 85
rect 9 83 10 85
rect 6 82 10 83
rect 18 85 22 86
rect 18 83 19 85
rect 21 83 22 85
rect 10 65 14 76
rect 10 63 11 65
rect 13 63 14 65
rect 10 45 14 63
rect 10 43 11 45
rect 13 43 14 45
rect 10 32 14 43
rect 18 46 22 83
rect 30 56 34 86
rect 28 55 34 56
rect 28 53 29 55
rect 31 53 34 55
rect 28 52 34 53
rect 18 45 24 46
rect 18 43 21 45
rect 23 43 24 45
rect 18 42 24 43
rect 18 27 22 42
rect 30 36 34 52
rect 28 35 34 36
rect 28 33 29 35
rect 31 33 34 35
rect 28 32 34 33
rect 6 25 22 27
rect 6 23 7 25
rect 9 23 22 25
rect 6 22 10 23
rect 30 22 34 32
rect 40 85 46 86
rect 40 83 43 85
rect 45 83 46 85
rect 40 82 46 83
rect 80 85 96 87
rect 80 83 81 85
rect 83 83 96 85
rect 80 82 84 83
rect 40 76 44 82
rect 40 75 46 76
rect 40 73 43 75
rect 45 73 46 75
rect 40 72 46 73
rect 40 66 44 72
rect 40 65 46 66
rect 40 63 43 65
rect 45 63 46 65
rect 40 62 46 63
rect 40 56 44 62
rect 40 52 48 56
rect 40 26 44 52
rect 84 45 88 76
rect 84 43 85 45
rect 87 43 88 45
rect 84 32 88 43
rect 92 46 96 83
rect 104 56 108 86
rect 102 55 108 56
rect 102 53 103 55
rect 105 53 108 55
rect 102 52 108 53
rect 92 45 98 46
rect 92 43 95 45
rect 97 43 98 45
rect 92 42 98 43
rect 40 25 46 26
rect 40 23 43 25
rect 45 23 46 25
rect 40 22 46 23
rect 92 25 96 42
rect 104 36 108 52
rect 102 35 108 36
rect 102 33 103 35
rect 105 33 108 35
rect 102 32 108 33
rect 92 23 93 25
rect 95 23 96 25
rect 92 22 96 23
rect 104 22 108 32
rect 114 85 120 86
rect 114 83 117 85
rect 119 83 120 85
rect 156 85 158 87
rect 160 85 198 87
rect 200 85 271 87
rect 273 85 302 87
rect 304 85 375 87
rect 377 85 397 87
rect 156 84 397 85
rect 429 85 433 92
rect 114 82 120 83
rect 114 76 118 82
rect 155 78 159 79
rect 114 75 120 76
rect 114 73 117 75
rect 119 73 120 75
rect 114 72 120 73
rect 155 74 168 78
rect 155 72 157 74
rect 114 66 118 72
rect 155 67 159 72
rect 114 65 120 66
rect 114 63 117 65
rect 119 63 120 65
rect 114 62 120 63
rect 155 65 157 67
rect 114 56 118 62
rect 114 52 122 56
rect 114 26 118 52
rect 155 46 159 65
rect 187 66 191 71
rect 187 64 188 66
rect 190 64 191 66
rect 187 62 191 64
rect 170 60 191 62
rect 170 58 184 60
rect 186 58 191 60
rect 195 70 200 72
rect 195 68 197 70
rect 199 68 200 70
rect 235 73 247 79
rect 195 66 200 68
rect 195 64 196 66
rect 198 64 200 66
rect 195 63 200 64
rect 195 61 197 63
rect 199 61 200 63
rect 195 59 200 61
rect 227 68 231 71
rect 227 66 228 68
rect 230 66 231 68
rect 155 44 160 46
rect 155 42 157 44
rect 159 42 160 44
rect 155 40 160 42
rect 170 53 191 54
rect 170 51 174 53
rect 176 51 188 53
rect 190 51 191 53
rect 170 50 191 51
rect 187 41 191 50
rect 195 39 199 59
rect 227 62 231 66
rect 218 61 231 62
rect 218 59 224 61
rect 226 59 231 61
rect 218 58 231 59
rect 235 68 240 73
rect 235 66 237 68
rect 239 66 240 68
rect 235 61 240 66
rect 235 59 237 61
rect 239 59 240 61
rect 235 57 240 59
rect 210 53 224 54
rect 210 51 214 53
rect 216 51 224 53
rect 210 50 224 51
rect 195 37 197 39
rect 199 37 207 39
rect 195 33 207 37
rect 219 44 224 50
rect 219 42 220 44
rect 222 42 224 44
rect 219 41 224 42
rect 251 48 256 55
rect 279 70 295 71
rect 279 68 281 70
rect 283 68 295 70
rect 279 66 295 68
rect 291 61 295 66
rect 291 59 292 61
rect 294 59 295 61
rect 251 47 253 48
rect 243 46 253 47
rect 255 46 256 48
rect 243 44 256 46
rect 243 42 245 44
rect 247 42 256 44
rect 243 41 256 42
rect 291 38 295 59
rect 271 37 295 38
rect 271 35 273 37
rect 275 35 295 37
rect 271 34 295 35
rect 299 70 304 72
rect 299 68 301 70
rect 303 68 304 70
rect 429 83 430 85
rect 432 83 433 85
rect 429 82 433 83
rect 441 85 489 86
rect 441 83 442 85
rect 444 83 486 85
rect 488 83 489 85
rect 441 82 489 83
rect 517 85 521 86
rect 517 83 518 85
rect 520 83 521 85
rect 339 73 351 79
rect 517 76 521 83
rect 541 85 545 86
rect 541 83 542 85
rect 544 83 545 85
rect 431 75 459 76
rect 299 63 304 68
rect 299 61 301 63
rect 303 61 304 63
rect 299 59 304 61
rect 331 68 335 71
rect 331 66 332 68
rect 334 66 335 68
rect 299 53 303 59
rect 299 51 300 53
rect 302 51 303 53
rect 299 39 303 51
rect 331 62 335 66
rect 322 61 335 62
rect 322 59 323 61
rect 325 59 328 61
rect 330 59 335 61
rect 322 58 335 59
rect 339 68 344 73
rect 339 66 341 68
rect 343 66 344 68
rect 339 61 344 66
rect 431 73 456 75
rect 458 73 459 75
rect 431 72 459 73
rect 465 75 534 76
rect 541 75 545 83
rect 465 73 466 75
rect 468 73 535 75
rect 465 72 535 73
rect 339 59 341 61
rect 343 59 344 61
rect 339 57 344 59
rect 314 53 328 54
rect 314 51 318 53
rect 320 51 328 53
rect 314 50 328 51
rect 299 37 301 39
rect 303 37 311 39
rect 299 33 311 37
rect 323 44 328 50
rect 323 42 324 44
rect 326 42 328 44
rect 323 41 328 42
rect 355 48 360 55
rect 383 70 399 71
rect 383 68 385 70
rect 387 68 399 70
rect 383 66 399 68
rect 355 47 357 48
rect 347 46 357 47
rect 359 46 360 48
rect 347 44 360 46
rect 347 42 349 44
rect 351 42 360 44
rect 347 41 360 42
rect 395 38 399 66
rect 431 56 435 72
rect 429 55 435 56
rect 429 53 430 55
rect 432 53 435 55
rect 429 52 435 53
rect 375 37 399 38
rect 375 35 377 37
rect 379 35 399 37
rect 375 34 399 35
rect 431 32 435 52
rect 441 65 473 66
rect 441 63 442 65
rect 444 63 470 65
rect 472 63 473 65
rect 441 62 473 63
rect 441 38 445 62
rect 451 55 455 56
rect 451 53 452 55
rect 454 53 455 55
rect 451 45 455 53
rect 462 55 475 56
rect 462 53 472 55
rect 474 53 475 55
rect 462 52 475 53
rect 481 46 485 72
rect 476 45 485 46
rect 475 43 485 45
rect 491 56 495 66
rect 501 65 511 66
rect 501 63 508 65
rect 510 63 511 65
rect 501 62 511 63
rect 517 65 524 66
rect 517 63 518 65
rect 520 63 525 65
rect 517 62 525 63
rect 507 56 511 62
rect 491 55 501 56
rect 491 53 498 55
rect 500 53 501 55
rect 491 52 501 53
rect 507 52 515 56
rect 475 42 484 43
rect 491 42 495 52
rect 507 46 511 52
rect 501 45 511 46
rect 501 43 508 45
rect 510 43 511 45
rect 501 42 511 43
rect 441 37 446 38
rect 441 35 442 37
rect 444 36 446 37
rect 475 36 479 42
rect 521 41 525 62
rect 518 40 525 41
rect 517 39 525 40
rect 517 37 518 39
rect 520 38 525 39
rect 520 37 524 38
rect 517 36 521 37
rect 444 35 459 36
rect 441 34 456 35
rect 442 33 456 34
rect 458 33 459 35
rect 442 32 459 33
rect 465 35 479 36
rect 465 33 466 35
rect 468 33 479 35
rect 487 35 521 36
rect 487 33 488 35
rect 490 33 504 35
rect 506 33 521 35
rect 465 32 478 33
rect 487 32 520 33
rect 156 27 399 28
rect 114 25 120 26
rect 114 23 117 25
rect 119 23 120 25
rect 114 22 120 23
rect 156 25 158 27
rect 160 25 198 27
rect 200 25 208 27
rect 210 25 238 27
rect 240 25 291 27
rect 293 25 302 27
rect 304 25 312 27
rect 314 25 342 27
rect 344 25 395 27
rect 397 25 399 27
rect 531 26 535 72
rect 541 73 542 75
rect 544 73 545 75
rect 541 65 545 73
rect 541 63 542 65
rect 544 63 545 65
rect 541 35 545 63
rect 553 85 557 92
rect 553 83 554 85
rect 556 83 557 85
rect 553 75 557 83
rect 553 73 554 75
rect 556 73 557 75
rect 553 65 557 73
rect 553 63 554 65
rect 556 63 557 65
rect 553 62 557 63
rect 565 75 569 76
rect 565 73 566 75
rect 568 73 569 75
rect 565 65 569 73
rect 565 63 566 65
rect 568 63 569 65
rect 541 33 542 35
rect 544 33 545 35
rect 541 32 545 33
rect 555 55 559 56
rect 555 53 556 55
rect 558 53 559 55
rect 555 37 559 53
rect 555 35 556 37
rect 558 35 559 37
rect 555 26 559 35
rect 156 16 399 25
rect 429 25 433 26
rect 429 23 430 25
rect 432 23 433 25
rect 429 16 433 23
rect 441 25 489 26
rect 441 23 442 25
rect 444 23 486 25
rect 488 23 489 25
rect 441 22 489 23
rect 517 25 559 26
rect 517 23 518 25
rect 520 23 559 25
rect 565 47 569 63
rect 565 45 566 47
rect 568 45 569 47
rect 565 27 569 45
rect 565 25 566 27
rect 568 25 569 27
rect 565 24 569 25
rect 517 22 558 23
rect 0 15 575 16
rect 0 13 31 15
rect 33 13 81 15
rect 83 13 105 15
rect 107 13 498 15
rect 500 13 530 15
rect 532 13 554 15
rect 556 13 575 15
rect 0 4 575 13
<< alu2 >>
rect 227 68 240 69
rect 187 66 200 68
rect 187 64 188 66
rect 190 64 196 66
rect 198 64 200 66
rect 227 66 228 68
rect 230 66 237 68
rect 239 66 240 68
rect 227 65 240 66
rect 331 68 344 69
rect 331 66 332 68
rect 334 66 341 68
rect 343 66 344 68
rect 331 65 344 66
rect 187 63 200 64
rect 291 61 326 62
rect 291 59 292 61
rect 294 59 323 61
rect 325 59 326 61
rect 291 58 326 59
rect 187 53 303 54
rect 187 51 188 53
rect 190 51 300 53
rect 302 51 303 53
rect 187 50 303 51
rect 219 44 251 46
rect 219 42 220 44
rect 222 42 245 44
rect 247 42 251 44
rect 219 41 251 42
rect 323 44 355 46
rect 323 42 324 44
rect 326 42 349 44
rect 351 42 355 44
rect 323 41 355 42
<< ptie >>
rect 156 27 162 29
rect 196 27 202 29
rect 156 25 158 27
rect 160 25 162 27
rect 156 23 162 25
rect 196 25 198 27
rect 200 25 202 27
rect 196 23 202 25
rect 236 27 242 29
rect 236 25 238 27
rect 240 25 242 27
rect 236 23 242 25
rect 300 27 306 29
rect 300 25 302 27
rect 304 25 306 27
rect 300 23 306 25
rect 340 27 346 29
rect 340 25 342 27
rect 344 25 346 27
rect 340 23 346 25
<< ntie >>
rect 79 99 97 101
rect 564 99 570 101
rect 79 97 81 99
rect 83 97 93 99
rect 95 97 97 99
rect 79 95 97 97
rect 156 87 162 89
rect 156 85 158 87
rect 160 85 162 87
rect 196 87 202 89
rect 156 83 162 85
rect 196 85 198 87
rect 200 85 202 87
rect 269 87 275 89
rect 196 83 202 85
rect 269 85 271 87
rect 273 85 275 87
rect 300 87 306 89
rect 269 83 275 85
rect 300 85 302 87
rect 304 85 306 87
rect 373 87 379 89
rect 300 83 306 85
rect 373 85 375 87
rect 377 85 379 87
rect 373 83 379 85
rect 564 97 566 99
rect 568 97 570 99
rect 564 89 570 97
<< nmos >>
rect 13 19 15 39
rect 162 37 164 46
rect 172 40 174 46
rect 182 40 184 46
rect 202 35 204 44
rect 25 9 27 29
rect 37 9 39 29
rect 87 19 89 29
rect 99 19 101 29
rect 111 9 113 29
rect 215 33 217 44
rect 222 33 224 44
rect 242 37 244 46
rect 258 32 260 41
rect 268 32 270 41
rect 278 29 280 41
rect 285 29 287 41
rect 306 35 308 44
rect 319 33 321 44
rect 326 33 328 44
rect 346 37 348 46
rect 362 32 364 41
rect 372 32 374 41
rect 382 29 384 41
rect 389 29 391 41
rect 436 33 438 41
rect 448 15 450 27
rect 460 15 462 27
rect 472 15 474 27
rect 480 15 482 27
rect 524 33 526 41
rect 492 11 494 23
rect 504 11 506 23
rect 512 11 514 23
rect 536 11 538 31
rect 548 11 550 31
rect 560 21 562 31
<< pmos >>
rect 13 69 15 89
rect 25 69 27 89
rect 37 59 39 99
rect 91 59 93 89
rect 99 59 101 89
rect 111 59 113 99
rect 162 58 164 76
rect 175 65 177 86
rect 182 65 184 86
rect 202 59 204 77
rect 212 66 214 79
rect 222 66 224 79
rect 250 59 252 86
rect 266 59 268 77
rect 276 59 278 77
rect 286 59 288 86
rect 306 59 308 77
rect 316 66 318 79
rect 326 66 328 79
rect 354 59 356 86
rect 370 59 372 77
rect 380 59 382 77
rect 390 59 392 86
rect 448 79 450 99
rect 460 79 462 99
rect 472 79 474 99
rect 480 79 482 99
rect 492 79 494 99
rect 504 79 506 99
rect 512 79 514 99
rect 436 59 438 73
rect 524 59 526 73
rect 536 59 538 99
rect 548 59 550 99
rect 560 59 562 79
<< polyct0 >>
rect 164 51 166 53
rect 204 51 206 53
rect 274 51 276 53
rect 284 52 286 54
rect 308 51 310 53
rect 378 51 380 53
rect 388 52 390 54
<< polyct1 >>
rect 11 63 13 65
rect 29 53 31 55
rect 11 43 13 45
rect 103 53 105 55
rect 21 43 23 45
rect 29 33 31 35
rect 85 43 87 45
rect 184 58 186 60
rect 174 51 176 53
rect 224 59 226 61
rect 237 59 239 61
rect 214 51 216 53
rect 95 43 97 45
rect 103 33 105 35
rect 328 59 330 61
rect 341 59 343 61
rect 253 46 255 48
rect 318 51 320 53
rect 430 53 432 55
rect 357 46 359 48
rect 456 73 458 75
rect 452 53 454 55
rect 470 63 472 65
rect 472 53 474 55
rect 456 33 458 35
rect 508 63 510 65
rect 498 53 500 55
rect 488 33 490 35
rect 508 43 510 45
rect 556 53 558 55
rect 566 45 568 47
rect 504 33 506 35
rect 556 35 558 37
<< ndifct0 >>
rect 177 42 179 44
rect 168 29 170 31
rect 237 42 239 44
rect 227 35 229 37
rect 251 34 253 36
rect 187 29 189 31
rect 263 37 265 39
rect 341 42 343 44
rect 331 35 333 37
rect 355 34 357 36
rect 367 37 369 39
<< ndifct1 >>
rect 7 23 9 25
rect 157 42 159 44
rect 197 37 199 39
rect 31 13 33 15
rect 43 23 45 25
rect 93 23 95 25
rect 81 13 83 15
rect 105 13 107 15
rect 117 23 119 25
rect 273 35 275 37
rect 208 25 210 27
rect 301 37 303 39
rect 291 25 293 27
rect 377 35 379 37
rect 312 25 314 27
rect 395 25 397 27
rect 442 35 444 37
rect 466 33 468 35
rect 430 23 432 25
rect 442 23 444 25
rect 486 23 488 25
rect 518 37 520 39
rect 542 33 544 35
rect 518 23 520 25
rect 498 13 500 15
rect 530 13 532 15
rect 566 25 568 27
rect 554 13 556 15
<< ntiect1 >>
rect 81 97 83 99
rect 93 97 95 99
rect 158 85 160 87
rect 198 85 200 87
rect 271 85 273 87
rect 302 85 304 87
rect 375 85 377 87
rect 566 97 568 99
<< ptiect1 >>
rect 158 25 160 27
rect 198 25 200 27
rect 238 25 240 27
rect 302 25 304 27
rect 342 25 344 27
<< pdifct0 >>
rect 168 82 170 84
rect 187 75 189 77
rect 207 73 209 75
rect 217 75 219 77
rect 217 68 219 70
rect 227 75 229 77
rect 245 61 247 63
rect 255 82 257 84
rect 255 75 257 77
rect 271 68 273 70
rect 271 61 273 63
rect 291 76 293 78
rect 311 73 313 75
rect 321 75 323 77
rect 321 68 323 70
rect 331 75 333 77
rect 349 61 351 63
rect 359 82 361 84
rect 359 75 361 77
rect 375 68 377 70
rect 375 61 377 63
rect 395 76 397 78
<< pdifct1 >>
rect 7 93 9 95
rect 31 93 33 95
rect 7 83 9 85
rect 19 83 21 85
rect 105 93 107 95
rect 43 83 45 85
rect 43 73 45 75
rect 43 63 45 65
rect 81 83 83 85
rect 117 83 119 85
rect 117 73 119 75
rect 117 63 119 65
rect 157 72 159 74
rect 157 65 159 67
rect 197 68 199 70
rect 197 61 199 63
rect 281 68 283 70
rect 301 68 303 70
rect 301 61 303 63
rect 385 68 387 70
rect 430 83 432 85
rect 442 83 444 85
rect 486 83 488 85
rect 498 93 500 95
rect 518 83 520 85
rect 530 95 532 97
rect 442 63 444 65
rect 466 73 468 75
rect 518 63 520 65
rect 542 83 544 85
rect 542 73 544 75
rect 542 63 544 65
rect 554 95 556 97
rect 554 83 556 85
rect 554 73 556 75
rect 554 63 556 65
rect 566 73 568 75
rect 566 63 568 65
<< alu0 >>
rect 166 82 168 84
rect 170 82 172 84
rect 166 81 172 82
rect 174 77 191 78
rect 174 75 187 77
rect 189 75 191 77
rect 174 74 191 75
rect 205 75 211 84
rect 159 63 160 74
rect 174 70 178 74
rect 205 73 207 75
rect 209 73 211 75
rect 205 72 211 73
rect 216 77 220 79
rect 216 75 217 77
rect 219 75 220 77
rect 163 66 178 70
rect 163 53 167 66
rect 216 70 220 75
rect 225 77 231 84
rect 254 82 255 84
rect 257 82 258 84
rect 225 75 227 77
rect 229 75 231 77
rect 225 74 231 75
rect 254 77 258 82
rect 254 75 255 77
rect 257 75 258 77
rect 254 73 258 75
rect 262 78 295 79
rect 262 76 291 78
rect 293 76 295 78
rect 262 75 295 76
rect 309 75 315 84
rect 216 69 217 70
rect 203 68 217 69
rect 219 68 220 70
rect 203 65 220 68
rect 182 57 188 58
rect 163 51 164 53
rect 166 51 167 53
rect 163 45 167 51
rect 163 44 181 45
rect 163 42 177 44
rect 179 42 181 44
rect 163 41 181 42
rect 203 53 207 65
rect 262 64 266 75
rect 309 73 311 75
rect 313 73 315 75
rect 309 72 315 73
rect 320 77 324 79
rect 320 75 321 77
rect 323 75 324 77
rect 243 63 266 64
rect 243 61 245 63
rect 247 61 266 63
rect 243 60 266 61
rect 243 54 247 60
rect 203 51 204 53
rect 206 51 207 53
rect 203 46 207 51
rect 203 42 215 46
rect 199 39 200 41
rect 211 38 215 42
rect 236 50 247 54
rect 236 44 240 50
rect 262 54 266 60
rect 270 70 274 72
rect 270 68 271 70
rect 273 68 274 70
rect 270 63 274 68
rect 270 61 271 63
rect 273 62 274 63
rect 273 61 286 62
rect 270 58 286 61
rect 282 56 286 58
rect 282 54 287 56
rect 262 53 278 54
rect 262 51 274 53
rect 276 51 278 53
rect 262 50 278 51
rect 282 52 284 54
rect 286 52 287 54
rect 282 50 287 52
rect 236 42 237 44
rect 239 42 240 44
rect 236 40 240 42
rect 282 46 286 50
rect 262 42 286 46
rect 262 39 266 42
rect 211 37 231 38
rect 262 37 263 39
rect 265 37 266 39
rect 211 35 227 37
rect 229 35 231 37
rect 211 34 231 35
rect 249 36 255 37
rect 249 34 251 36
rect 253 34 255 36
rect 262 35 266 37
rect 320 70 324 75
rect 329 77 335 84
rect 358 82 359 84
rect 361 82 362 84
rect 329 75 331 77
rect 333 75 335 77
rect 329 74 335 75
rect 358 77 362 82
rect 358 75 359 77
rect 361 75 362 77
rect 358 73 362 75
rect 366 78 399 79
rect 366 76 395 78
rect 397 76 399 78
rect 366 75 399 76
rect 320 69 321 70
rect 307 68 321 69
rect 323 68 324 70
rect 307 65 324 68
rect 307 53 311 65
rect 366 64 370 75
rect 347 63 370 64
rect 347 61 349 63
rect 351 61 370 63
rect 347 60 370 61
rect 347 54 351 60
rect 307 51 308 53
rect 310 51 311 53
rect 307 46 311 51
rect 307 42 319 46
rect 303 39 304 41
rect 166 31 172 32
rect 166 29 168 31
rect 170 29 172 31
rect 166 28 172 29
rect 185 31 191 32
rect 185 29 187 31
rect 189 29 191 31
rect 185 28 191 29
rect 249 28 255 34
rect 315 38 319 42
rect 340 50 351 54
rect 340 44 344 50
rect 366 54 370 60
rect 374 70 378 72
rect 374 68 375 70
rect 377 68 378 70
rect 374 63 378 68
rect 374 61 375 63
rect 377 62 378 63
rect 377 61 390 62
rect 374 58 390 61
rect 386 56 390 58
rect 386 54 391 56
rect 366 53 382 54
rect 366 51 378 53
rect 380 51 382 53
rect 366 50 382 51
rect 386 52 388 54
rect 390 52 391 54
rect 386 50 391 52
rect 340 42 341 44
rect 343 42 344 44
rect 340 40 344 42
rect 386 46 390 50
rect 366 42 390 46
rect 366 39 370 42
rect 315 37 335 38
rect 366 37 367 39
rect 369 37 370 39
rect 315 35 331 37
rect 333 35 335 37
rect 315 34 335 35
rect 353 36 359 37
rect 353 34 355 36
rect 357 34 359 36
rect 366 35 370 37
rect 353 28 359 34
<< via1 >>
rect 188 64 190 66
rect 196 64 198 66
rect 228 66 230 68
rect 188 51 190 53
rect 237 66 239 68
rect 220 42 222 44
rect 292 59 294 61
rect 245 42 247 44
rect 332 66 334 68
rect 300 51 302 53
rect 323 59 325 61
rect 341 66 343 68
rect 324 42 326 44
rect 349 42 351 44
<< labels >>
rlabel alu1 12 54 12 54 6 i0
rlabel alu1 27 10 27 10 6 vss
rlabel alu1 32 54 32 54 6 i1
rlabel alu1 27 98 27 98 6 vdd
rlabel alu1 86 54 86 54 6 i1
rlabel alu1 101 10 101 10 6 vss
rlabel alu1 106 54 106 54 6 i0
rlabel alu1 101 98 101 98 6 vdd
rlabel alu0 238 47 238 47 6 bn
rlabel alu0 284 52 284 52 6 an
rlabel alu1 265 24 265 24 6 vss
rlabel alu1 265 88 265 88 6 vdd
rlabel alu1 213 88 213 88 6 vdd
rlabel alu1 213 24 213 24 6 vss
rlabel alu0 205 55 205 55 6 zn
rlabel alu1 317 24 317 24 6 vss
rlabel alu1 317 88 317 88 6 vdd
rlabel alu1 397 48 397 48 1 sum
rlabel alu1 369 88 369 88 6 vdd
rlabel alu1 369 24 369 24 6 vss
rlabel alu1 293 48 293 48 1 s
rlabel alu1 317 51 317 51 1 cin
rlabel alu1 205 36 205 36 1 co
rlabel alu0 309 54 309 54 1 zn_1
rlabel alu0 342 47 342 47 1 bn_1
rlabel alu0 368 39 368 39 1 an_1
rlabel alu1 173 88 173 88 6 vdd
rlabel alu1 173 24 173 24 6 vss
rlabel alu1 309 36 309 36 1 c1
rlabel alu1 157 56 157 56 1 cout
rlabel alu0 182 76 182 76 1 zn_2
rlabel alu1 433 54 433 54 6 cmd1
rlabel polyct1 453 54 453 54 6 i2
rlabel polyct1 473 54 473 54 6 i1
rlabel alu1 498 10 498 10 6 vss
rlabel alu1 503 44 503 44 6 i0
rlabel alu1 493 54 493 54 6 cmd0
rlabel alu1 503 64 503 64 6 i0
rlabel alu1 498 98 498 98 6 vdd
rlabel alu1 513 54 513 54 6 i0
rlabel alu1 543 59 543 59 6 nq
rlabel alu1 42 54 42 54 1 andout
rlabel alu1 116 54 116 54 1 orout
rlabel alu2 213 52 213 52 1 in1
rlabel via1 229 67 229 67 1 in2
rlabel polyct1 253 48 253 48 1 in1
<< end >>
