magic
tech scmos
timestamp 1608962259
<< ab >>
rect 68 581 74 586
rect 172 581 178 586
rect 5 573 654 581
rect 5 549 253 573
rect 5 517 68 549
rect 69 536 172 549
rect 173 545 253 549
rect 254 545 654 573
rect 173 536 654 545
rect 69 523 654 536
rect 69 517 172 523
rect 173 517 253 523
rect 254 517 654 523
rect 5 514 654 517
rect 3 511 654 514
rect 3 508 11 511
rect 253 508 654 511
rect 5 501 654 508
rect 5 469 85 501
rect 86 469 189 501
rect 190 495 253 501
rect 254 495 654 501
rect 190 483 654 495
rect 190 469 253 483
rect 5 445 253 469
rect 254 445 654 483
rect 5 439 654 445
rect 3 437 654 439
rect 5 429 654 437
rect 5 405 253 429
rect 5 373 68 405
rect 69 392 172 405
rect 173 392 253 405
rect 69 390 253 392
rect 254 390 654 429
rect 69 380 654 390
rect 69 373 172 380
rect 173 373 253 380
rect 254 373 654 380
rect 5 371 654 373
rect 3 363 654 371
rect 5 357 654 363
rect 5 325 85 357
rect 86 325 189 357
rect 190 344 253 357
rect 254 344 654 357
rect 190 339 654 344
rect 190 325 253 339
rect 5 319 253 325
rect 254 319 654 339
rect 5 314 654 319
rect 5 301 253 314
rect 254 301 654 314
rect 5 285 654 301
rect 5 261 253 285
rect 5 229 68 261
rect 69 248 172 261
rect 173 257 253 261
rect 254 257 654 285
rect 173 248 654 257
rect 69 235 654 248
rect 69 229 172 235
rect 173 229 253 235
rect 254 229 654 235
rect 5 226 654 229
rect 3 223 654 226
rect 3 220 11 223
rect 253 220 654 223
rect 5 213 654 220
rect 5 181 85 213
rect 86 181 189 213
rect 190 207 253 213
rect 254 207 654 213
rect 190 195 654 207
rect 190 181 253 195
rect 5 157 253 181
rect 254 157 654 195
rect 5 151 654 157
rect 3 149 654 151
rect 5 141 654 149
rect 5 117 253 141
rect 5 85 68 117
rect 69 104 172 117
rect 173 104 253 117
rect 69 92 253 104
rect 69 85 172 92
rect 173 85 253 92
rect 254 85 654 141
rect 5 83 654 85
rect 3 75 654 83
rect 5 69 654 75
rect 5 37 85 69
rect 86 37 189 69
rect 190 56 253 69
rect 254 56 654 69
rect 190 51 654 56
rect 190 37 253 51
rect 5 31 253 37
rect 254 31 654 51
rect 5 26 654 31
rect 5 13 253 26
rect 254 13 654 26
rect 5 5 654 13
rect 80 0 86 5
rect 184 0 190 5
<< nwell >>
rect 0 469 659 549
rect 0 325 659 405
rect 0 181 659 261
rect 0 37 659 117
<< pwell >>
rect 0 549 659 586
rect 0 405 659 469
rect 0 261 659 325
rect 0 117 659 181
rect 0 0 659 37
<< poly >>
rect 32 577 57 579
rect 15 572 17 577
rect 22 572 24 577
rect 32 569 34 577
rect 42 569 44 573
rect 55 569 57 577
rect 55 567 60 569
rect 78 568 80 573
rect 85 568 87 573
rect 136 577 161 579
rect 119 572 121 577
rect 126 572 128 577
rect 58 564 60 567
rect 15 551 17 560
rect 22 557 24 560
rect 22 555 26 557
rect 32 556 34 560
rect 42 557 44 560
rect 24 552 26 555
rect 42 555 51 557
rect 98 566 100 570
rect 136 569 138 577
rect 146 569 148 573
rect 159 569 161 577
rect 159 567 164 569
rect 182 568 184 573
rect 189 568 191 573
rect 162 564 164 567
rect 42 553 47 555
rect 49 553 51 555
rect 14 549 20 551
rect 14 547 16 549
rect 18 547 20 549
rect 14 545 20 547
rect 24 550 30 552
rect 24 548 26 550
rect 28 548 30 550
rect 24 546 30 548
rect 42 551 51 553
rect 42 547 44 551
rect 58 547 60 555
rect 14 542 16 545
rect 24 542 26 546
rect 34 545 44 547
rect 50 545 63 547
rect 34 542 36 545
rect 50 542 52 545
rect 61 544 63 545
rect 78 544 80 557
rect 85 552 87 557
rect 98 552 100 557
rect 84 550 90 552
rect 84 548 86 550
rect 88 548 90 550
rect 84 546 90 548
rect 94 550 100 552
rect 119 551 121 560
rect 126 557 128 560
rect 126 555 130 557
rect 136 556 138 560
rect 146 557 148 560
rect 128 552 130 555
rect 146 555 155 557
rect 202 566 204 570
rect 281 577 306 579
rect 264 572 266 577
rect 271 572 273 577
rect 222 561 224 566
rect 232 561 234 566
rect 242 564 244 569
rect 146 553 151 555
rect 153 553 155 555
rect 94 548 96 550
rect 98 548 100 550
rect 94 546 100 548
rect 61 542 67 544
rect 24 520 26 524
rect 34 520 36 524
rect 14 511 16 515
rect 61 540 63 542
rect 65 540 67 542
rect 61 538 67 540
rect 74 542 80 544
rect 74 540 76 542
rect 78 540 80 542
rect 74 538 80 540
rect 78 535 80 538
rect 88 535 90 546
rect 98 542 100 546
rect 118 549 124 551
rect 118 547 120 549
rect 122 547 124 549
rect 118 545 124 547
rect 128 550 134 552
rect 128 548 130 550
rect 132 548 134 550
rect 128 546 134 548
rect 146 551 155 553
rect 146 547 148 551
rect 162 547 164 555
rect 118 542 120 545
rect 128 542 130 546
rect 138 545 148 547
rect 154 545 167 547
rect 138 542 140 545
rect 154 542 156 545
rect 165 544 167 545
rect 182 544 184 557
rect 189 552 191 557
rect 202 552 204 557
rect 281 569 283 577
rect 291 569 293 573
rect 304 569 306 577
rect 304 567 309 569
rect 327 568 329 573
rect 334 568 336 573
rect 307 564 309 567
rect 188 550 194 552
rect 188 548 190 550
rect 192 548 194 550
rect 188 546 194 548
rect 198 550 204 552
rect 198 548 200 550
rect 202 548 204 550
rect 198 546 204 548
rect 165 542 171 544
rect 78 517 80 522
rect 88 517 90 522
rect 98 520 100 524
rect 50 511 52 515
rect 128 520 130 524
rect 138 520 140 524
rect 118 511 120 515
rect 165 540 167 542
rect 169 540 171 542
rect 165 538 171 540
rect 178 542 184 544
rect 178 540 180 542
rect 182 540 184 542
rect 178 538 184 540
rect 182 535 184 538
rect 192 535 194 546
rect 202 542 204 546
rect 222 545 224 555
rect 232 552 234 555
rect 242 552 244 555
rect 228 550 234 552
rect 228 548 230 550
rect 232 548 234 550
rect 228 546 234 548
rect 238 550 244 552
rect 264 551 266 560
rect 271 557 273 560
rect 271 555 275 557
rect 281 556 283 560
rect 291 557 293 560
rect 273 552 275 555
rect 291 555 300 557
rect 347 566 349 570
rect 410 577 435 579
rect 410 569 412 577
rect 423 569 425 573
rect 433 569 435 577
rect 443 572 445 577
rect 450 572 452 577
rect 367 561 369 566
rect 377 561 379 566
rect 387 564 389 569
rect 407 567 412 569
rect 407 564 409 567
rect 291 553 296 555
rect 298 553 300 555
rect 238 548 240 550
rect 242 548 244 550
rect 238 546 244 548
rect 218 543 224 545
rect 218 541 220 543
rect 222 541 224 543
rect 218 539 224 541
rect 222 536 224 539
rect 229 536 231 546
rect 242 543 244 546
rect 263 549 269 551
rect 263 547 265 549
rect 267 547 269 549
rect 263 545 269 547
rect 273 550 279 552
rect 273 548 275 550
rect 277 548 279 550
rect 273 546 279 548
rect 291 551 300 553
rect 291 547 293 551
rect 307 547 309 555
rect 182 517 184 522
rect 192 517 194 522
rect 202 520 204 524
rect 154 511 156 515
rect 263 542 265 545
rect 273 542 275 546
rect 283 545 293 547
rect 299 545 312 547
rect 283 542 285 545
rect 299 542 301 545
rect 310 544 312 545
rect 327 544 329 557
rect 334 552 336 557
rect 347 552 349 557
rect 471 577 490 579
rect 471 567 473 577
rect 481 569 483 573
rect 488 569 490 577
rect 535 577 554 579
rect 498 569 500 574
rect 505 569 507 574
rect 515 569 517 574
rect 423 557 425 560
rect 416 555 425 557
rect 433 556 435 560
rect 443 557 445 560
rect 333 550 339 552
rect 333 548 335 550
rect 337 548 339 550
rect 333 546 339 548
rect 343 550 349 552
rect 343 548 345 550
rect 347 548 349 550
rect 343 546 349 548
rect 310 542 316 544
rect 242 520 244 525
rect 222 511 224 515
rect 229 511 231 515
rect 273 520 275 524
rect 283 520 285 524
rect 263 511 265 515
rect 310 540 312 542
rect 314 540 316 542
rect 310 538 316 540
rect 323 542 329 544
rect 323 540 325 542
rect 327 540 329 542
rect 323 538 329 540
rect 327 535 329 538
rect 337 535 339 546
rect 347 542 349 546
rect 367 545 369 555
rect 377 552 379 555
rect 387 552 389 555
rect 373 550 379 552
rect 373 548 375 550
rect 377 548 379 550
rect 373 546 379 548
rect 383 550 389 552
rect 383 548 385 550
rect 387 548 389 550
rect 383 546 389 548
rect 407 547 409 555
rect 416 553 418 555
rect 420 553 425 555
rect 416 551 425 553
rect 441 555 445 557
rect 441 552 443 555
rect 423 547 425 551
rect 437 550 443 552
rect 450 551 452 560
rect 437 548 439 550
rect 441 548 443 550
rect 363 543 369 545
rect 363 541 365 543
rect 367 541 369 543
rect 363 539 369 541
rect 367 536 369 539
rect 374 536 376 546
rect 387 543 389 546
rect 404 545 417 547
rect 423 545 433 547
rect 437 546 443 548
rect 404 544 406 545
rect 327 517 329 522
rect 337 517 339 522
rect 347 520 349 524
rect 299 511 301 515
rect 400 542 406 544
rect 415 542 417 545
rect 431 542 433 545
rect 441 542 443 546
rect 447 549 453 551
rect 447 547 449 549
rect 451 547 453 549
rect 447 545 453 547
rect 451 542 453 545
rect 471 543 473 561
rect 481 552 483 561
rect 477 550 483 552
rect 477 548 479 550
rect 481 548 483 550
rect 477 546 483 548
rect 488 548 490 561
rect 498 558 500 561
rect 494 556 500 558
rect 494 554 496 556
rect 498 554 500 556
rect 494 552 500 554
rect 488 546 500 548
rect 505 547 507 561
rect 535 567 537 577
rect 545 569 547 573
rect 552 569 554 577
rect 599 577 618 579
rect 562 569 564 574
rect 569 569 571 574
rect 579 569 581 574
rect 515 557 517 560
rect 512 555 518 557
rect 512 553 514 555
rect 516 553 518 555
rect 512 551 518 553
rect 400 540 402 542
rect 404 540 406 542
rect 400 538 406 540
rect 387 520 389 525
rect 367 511 369 515
rect 374 511 376 515
rect 431 520 433 524
rect 441 520 443 524
rect 415 511 417 515
rect 471 532 473 535
rect 464 530 473 532
rect 481 531 483 546
rect 487 540 493 542
rect 487 538 489 540
rect 491 538 493 540
rect 487 536 493 538
rect 488 531 490 536
rect 498 531 500 546
rect 504 545 510 547
rect 504 543 506 545
rect 508 543 510 545
rect 504 541 510 543
rect 505 531 507 541
rect 515 533 517 551
rect 535 543 537 561
rect 545 552 547 561
rect 541 550 547 552
rect 541 548 543 550
rect 545 548 547 550
rect 541 546 547 548
rect 552 548 554 561
rect 562 558 564 561
rect 558 556 564 558
rect 558 554 560 556
rect 562 554 564 556
rect 558 552 564 554
rect 552 546 564 548
rect 569 547 571 561
rect 599 567 601 577
rect 609 569 611 573
rect 616 569 618 577
rect 626 569 628 574
rect 633 569 635 574
rect 643 569 645 574
rect 579 557 581 560
rect 576 555 582 557
rect 576 553 578 555
rect 580 553 582 555
rect 576 551 582 553
rect 464 528 466 530
rect 468 528 470 530
rect 464 526 470 528
rect 535 532 537 535
rect 528 530 537 532
rect 545 531 547 546
rect 551 540 557 542
rect 551 538 553 540
rect 555 538 557 540
rect 551 536 557 538
rect 552 531 554 536
rect 562 531 564 546
rect 568 545 574 547
rect 568 543 570 545
rect 572 543 574 545
rect 568 541 574 543
rect 569 531 571 541
rect 579 533 581 551
rect 599 543 601 561
rect 609 552 611 561
rect 605 550 611 552
rect 605 548 607 550
rect 609 548 611 550
rect 605 546 611 548
rect 616 548 618 561
rect 626 558 628 561
rect 622 556 628 558
rect 622 554 624 556
rect 626 554 628 556
rect 622 552 628 554
rect 616 546 628 548
rect 633 547 635 561
rect 643 557 645 560
rect 640 555 646 557
rect 640 553 642 555
rect 644 553 646 555
rect 640 551 646 553
rect 528 528 530 530
rect 532 528 534 530
rect 528 526 534 528
rect 599 532 601 535
rect 592 530 601 532
rect 609 531 611 546
rect 615 540 621 542
rect 615 538 617 540
rect 619 538 621 540
rect 615 536 621 538
rect 616 531 618 536
rect 626 531 628 546
rect 632 545 638 547
rect 632 543 634 545
rect 636 543 638 545
rect 632 541 638 543
rect 633 531 635 541
rect 643 533 645 551
rect 592 528 594 530
rect 596 528 598 530
rect 592 526 598 528
rect 451 511 453 515
rect 481 511 483 515
rect 488 511 490 515
rect 498 511 500 515
rect 505 511 507 515
rect 515 511 517 515
rect 545 511 547 515
rect 552 511 554 515
rect 562 511 564 515
rect 569 511 571 515
rect 579 511 581 515
rect 609 511 611 515
rect 616 511 618 515
rect 626 511 628 515
rect 633 511 635 515
rect 643 511 645 515
rect 27 503 29 507
rect 34 503 36 507
rect 14 493 16 498
rect 102 503 104 507
rect 54 494 56 498
rect 64 496 66 501
rect 74 496 76 501
rect 14 472 16 475
rect 27 472 29 482
rect 34 479 36 482
rect 34 477 40 479
rect 34 475 36 477
rect 38 475 40 477
rect 34 473 40 475
rect 14 470 20 472
rect 14 468 16 470
rect 18 468 20 470
rect 14 466 20 468
rect 24 470 30 472
rect 24 468 26 470
rect 28 468 30 470
rect 24 466 30 468
rect 14 463 16 466
rect 24 463 26 466
rect 34 463 36 473
rect 54 472 56 476
rect 64 472 66 483
rect 74 480 76 483
rect 74 478 80 480
rect 74 476 76 478
rect 78 476 80 478
rect 74 474 80 476
rect 87 478 93 480
rect 87 476 89 478
rect 91 476 93 478
rect 138 503 140 507
rect 118 494 120 498
rect 128 494 130 498
rect 206 503 208 507
rect 158 494 160 498
rect 168 496 170 501
rect 178 496 180 501
rect 87 474 93 476
rect 54 470 60 472
rect 54 468 56 470
rect 58 468 60 470
rect 54 466 60 468
rect 64 470 70 472
rect 64 468 66 470
rect 68 468 70 470
rect 64 466 70 468
rect 54 461 56 466
rect 67 461 69 466
rect 74 461 76 474
rect 91 473 93 474
rect 102 473 104 476
rect 118 473 120 476
rect 91 471 104 473
rect 110 471 120 473
rect 128 472 130 476
rect 138 473 140 476
rect 94 463 96 471
rect 110 467 112 471
rect 103 465 112 467
rect 124 470 130 472
rect 124 468 126 470
rect 128 468 130 470
rect 124 466 130 468
rect 134 471 140 473
rect 134 469 136 471
rect 138 469 140 471
rect 134 467 140 469
rect 158 472 160 476
rect 168 472 170 483
rect 178 480 180 483
rect 178 478 184 480
rect 178 476 180 478
rect 182 476 184 478
rect 178 474 184 476
rect 191 478 197 480
rect 191 476 193 478
rect 195 476 197 478
rect 242 503 244 507
rect 263 503 265 507
rect 222 494 224 498
rect 232 494 234 498
rect 299 503 301 507
rect 273 494 275 498
rect 283 494 285 498
rect 367 503 369 507
rect 374 503 376 507
rect 327 496 329 501
rect 337 496 339 501
rect 347 494 349 498
rect 327 480 329 483
rect 310 478 316 480
rect 310 476 312 478
rect 314 476 316 478
rect 191 474 197 476
rect 158 470 164 472
rect 158 468 160 470
rect 162 468 164 470
rect 103 463 105 465
rect 107 463 112 465
rect 14 449 16 454
rect 24 452 26 457
rect 34 452 36 457
rect 54 448 56 452
rect 103 461 112 463
rect 128 463 130 466
rect 110 458 112 461
rect 120 458 122 462
rect 128 461 132 463
rect 130 458 132 461
rect 137 458 139 467
rect 158 466 164 468
rect 168 470 174 472
rect 168 468 170 470
rect 172 468 174 470
rect 168 466 174 468
rect 158 461 160 466
rect 171 461 173 466
rect 178 461 180 474
rect 195 473 197 474
rect 206 473 208 476
rect 222 473 224 476
rect 195 471 208 473
rect 214 471 224 473
rect 232 472 234 476
rect 242 473 244 476
rect 198 463 200 471
rect 214 467 216 471
rect 207 465 216 467
rect 228 470 234 472
rect 228 468 230 470
rect 232 468 234 470
rect 228 466 234 468
rect 238 471 244 473
rect 238 469 240 471
rect 242 469 244 471
rect 238 467 244 469
rect 263 473 265 476
rect 263 471 269 473
rect 263 469 265 471
rect 267 469 269 471
rect 263 467 269 469
rect 273 472 275 476
rect 283 473 285 476
rect 299 473 301 476
rect 310 474 316 476
rect 323 478 329 480
rect 323 476 325 478
rect 327 476 329 478
rect 323 474 329 476
rect 310 473 312 474
rect 273 470 279 472
rect 283 471 293 473
rect 299 471 312 473
rect 273 468 275 470
rect 277 468 279 470
rect 207 463 209 465
rect 211 463 216 465
rect 94 451 96 454
rect 67 445 69 450
rect 74 445 76 450
rect 94 449 99 451
rect 97 441 99 449
rect 110 445 112 449
rect 120 441 122 449
rect 158 448 160 452
rect 207 461 216 463
rect 232 463 234 466
rect 214 458 216 461
rect 224 458 226 462
rect 232 461 236 463
rect 234 458 236 461
rect 241 458 243 467
rect 264 458 266 467
rect 273 466 279 468
rect 291 467 293 471
rect 273 463 275 466
rect 271 461 275 463
rect 291 465 300 467
rect 291 463 296 465
rect 298 463 300 465
rect 307 463 309 471
rect 271 458 273 461
rect 281 458 283 462
rect 291 461 300 463
rect 291 458 293 461
rect 198 451 200 454
rect 130 441 132 446
rect 137 441 139 446
rect 97 439 122 441
rect 171 445 173 450
rect 178 445 180 450
rect 198 449 203 451
rect 201 441 203 449
rect 214 445 216 449
rect 224 441 226 449
rect 234 441 236 446
rect 241 441 243 446
rect 201 439 226 441
rect 327 461 329 474
rect 337 472 339 483
rect 415 503 417 507
rect 387 493 389 498
rect 367 479 369 482
rect 363 477 369 479
rect 347 472 349 476
rect 363 475 365 477
rect 367 475 369 477
rect 363 473 369 475
rect 333 470 339 472
rect 333 468 335 470
rect 337 468 339 470
rect 333 466 339 468
rect 343 470 349 472
rect 343 468 345 470
rect 347 468 349 470
rect 343 466 349 468
rect 334 461 336 466
rect 347 461 349 466
rect 367 463 369 473
rect 374 472 376 482
rect 400 478 406 480
rect 400 476 402 478
rect 404 476 406 478
rect 451 503 453 507
rect 481 503 483 507
rect 488 503 490 507
rect 498 503 500 507
rect 505 503 507 507
rect 515 503 517 507
rect 545 503 547 507
rect 552 503 554 507
rect 562 503 564 507
rect 569 503 571 507
rect 579 503 581 507
rect 609 503 611 507
rect 616 503 618 507
rect 626 503 628 507
rect 633 503 635 507
rect 643 503 645 507
rect 431 494 433 498
rect 441 494 443 498
rect 464 490 470 492
rect 464 488 466 490
rect 468 488 470 490
rect 464 486 473 488
rect 471 483 473 486
rect 387 472 389 475
rect 400 474 406 476
rect 373 470 379 472
rect 373 468 375 470
rect 377 468 379 470
rect 373 466 379 468
rect 383 470 389 472
rect 404 473 406 474
rect 415 473 417 476
rect 431 473 433 476
rect 404 471 417 473
rect 423 471 433 473
rect 441 472 443 476
rect 451 473 453 476
rect 383 468 385 470
rect 387 468 389 470
rect 383 466 389 468
rect 377 463 379 466
rect 387 463 389 466
rect 407 463 409 471
rect 423 467 425 471
rect 416 465 425 467
rect 437 470 443 472
rect 437 468 439 470
rect 441 468 443 470
rect 437 466 443 468
rect 447 471 453 473
rect 447 469 449 471
rect 451 469 453 471
rect 447 467 453 469
rect 416 463 418 465
rect 420 463 425 465
rect 307 451 309 454
rect 304 449 309 451
rect 264 441 266 446
rect 271 441 273 446
rect 281 441 283 449
rect 291 445 293 449
rect 304 441 306 449
rect 281 439 306 441
rect 327 445 329 450
rect 334 445 336 450
rect 347 448 349 452
rect 367 452 369 457
rect 377 452 379 457
rect 416 461 425 463
rect 441 463 443 466
rect 423 458 425 461
rect 433 458 435 462
rect 441 461 445 463
rect 443 458 445 461
rect 450 458 452 467
rect 387 449 389 454
rect 407 451 409 454
rect 407 449 412 451
rect 410 441 412 449
rect 423 445 425 449
rect 433 441 435 449
rect 471 457 473 475
rect 481 472 483 487
rect 488 482 490 487
rect 487 480 493 482
rect 487 478 489 480
rect 491 478 493 480
rect 487 476 493 478
rect 498 472 500 487
rect 505 477 507 487
rect 528 490 534 492
rect 528 488 530 490
rect 532 488 534 490
rect 528 486 537 488
rect 477 470 483 472
rect 477 468 479 470
rect 481 468 483 470
rect 477 466 483 468
rect 481 457 483 466
rect 488 470 500 472
rect 504 475 510 477
rect 504 473 506 475
rect 508 473 510 475
rect 504 471 510 473
rect 488 457 490 470
rect 494 464 500 466
rect 494 462 496 464
rect 498 462 500 464
rect 494 460 500 462
rect 498 457 500 460
rect 505 457 507 471
rect 515 467 517 485
rect 535 483 537 486
rect 512 465 518 467
rect 512 463 514 465
rect 516 463 518 465
rect 512 461 518 463
rect 515 458 517 461
rect 443 441 445 446
rect 450 441 452 446
rect 410 439 435 441
rect 471 441 473 451
rect 535 457 537 475
rect 545 472 547 487
rect 552 482 554 487
rect 551 480 557 482
rect 551 478 553 480
rect 555 478 557 480
rect 551 476 557 478
rect 562 472 564 487
rect 569 477 571 487
rect 592 490 598 492
rect 592 488 594 490
rect 596 488 598 490
rect 592 486 601 488
rect 541 470 547 472
rect 541 468 543 470
rect 545 468 547 470
rect 541 466 547 468
rect 545 457 547 466
rect 552 470 564 472
rect 568 475 574 477
rect 568 473 570 475
rect 572 473 574 475
rect 568 471 574 473
rect 552 457 554 470
rect 558 464 564 466
rect 558 462 560 464
rect 562 462 564 464
rect 558 460 564 462
rect 562 457 564 460
rect 569 457 571 471
rect 579 467 581 485
rect 599 483 601 486
rect 576 465 582 467
rect 576 463 578 465
rect 580 463 582 465
rect 576 461 582 463
rect 579 458 581 461
rect 481 445 483 449
rect 488 441 490 449
rect 498 444 500 449
rect 505 444 507 449
rect 515 444 517 449
rect 471 439 490 441
rect 535 441 537 451
rect 599 457 601 475
rect 609 472 611 487
rect 616 482 618 487
rect 615 480 621 482
rect 615 478 617 480
rect 619 478 621 480
rect 615 476 621 478
rect 626 472 628 487
rect 633 477 635 487
rect 605 470 611 472
rect 605 468 607 470
rect 609 468 611 470
rect 605 466 611 468
rect 609 457 611 466
rect 616 470 628 472
rect 632 475 638 477
rect 632 473 634 475
rect 636 473 638 475
rect 632 471 638 473
rect 616 457 618 470
rect 622 464 628 466
rect 622 462 624 464
rect 626 462 628 464
rect 622 460 628 462
rect 626 457 628 460
rect 633 457 635 471
rect 643 467 645 485
rect 640 465 646 467
rect 640 463 642 465
rect 644 463 646 465
rect 640 461 646 463
rect 643 458 645 461
rect 545 445 547 449
rect 552 441 554 449
rect 562 444 564 449
rect 569 444 571 449
rect 579 444 581 449
rect 535 439 554 441
rect 599 441 601 451
rect 609 445 611 449
rect 616 441 618 449
rect 626 444 628 449
rect 633 444 635 449
rect 643 444 645 449
rect 599 439 618 441
rect 32 433 57 435
rect 15 428 17 433
rect 22 428 24 433
rect 32 425 34 433
rect 42 425 44 429
rect 55 425 57 433
rect 55 423 60 425
rect 78 424 80 429
rect 85 424 87 429
rect 136 433 161 435
rect 119 428 121 433
rect 126 428 128 433
rect 58 420 60 423
rect 15 407 17 416
rect 22 413 24 416
rect 22 411 26 413
rect 32 412 34 416
rect 42 413 44 416
rect 24 408 26 411
rect 42 411 51 413
rect 98 422 100 426
rect 136 425 138 433
rect 146 425 148 429
rect 159 425 161 433
rect 159 423 164 425
rect 182 424 184 429
rect 189 424 191 429
rect 162 420 164 423
rect 42 409 47 411
rect 49 409 51 411
rect 14 405 20 407
rect 14 403 16 405
rect 18 403 20 405
rect 14 401 20 403
rect 24 406 30 408
rect 24 404 26 406
rect 28 404 30 406
rect 24 402 30 404
rect 42 407 51 409
rect 42 403 44 407
rect 58 403 60 411
rect 14 398 16 401
rect 24 398 26 402
rect 34 401 44 403
rect 50 401 63 403
rect 34 398 36 401
rect 50 398 52 401
rect 61 400 63 401
rect 78 400 80 413
rect 85 408 87 413
rect 98 408 100 413
rect 84 406 90 408
rect 84 404 86 406
rect 88 404 90 406
rect 84 402 90 404
rect 94 406 100 408
rect 119 407 121 416
rect 126 413 128 416
rect 126 411 130 413
rect 136 412 138 416
rect 146 413 148 416
rect 128 408 130 411
rect 146 411 155 413
rect 202 422 204 426
rect 281 433 306 435
rect 264 428 266 433
rect 271 428 273 433
rect 222 417 224 422
rect 232 417 234 422
rect 242 420 244 425
rect 146 409 151 411
rect 153 409 155 411
rect 94 404 96 406
rect 98 404 100 406
rect 94 402 100 404
rect 61 398 67 400
rect 24 376 26 380
rect 34 376 36 380
rect 14 367 16 371
rect 61 396 63 398
rect 65 396 67 398
rect 61 394 67 396
rect 74 398 80 400
rect 74 396 76 398
rect 78 396 80 398
rect 74 394 80 396
rect 78 391 80 394
rect 88 391 90 402
rect 98 398 100 402
rect 118 405 124 407
rect 118 403 120 405
rect 122 403 124 405
rect 118 401 124 403
rect 128 406 134 408
rect 128 404 130 406
rect 132 404 134 406
rect 128 402 134 404
rect 146 407 155 409
rect 146 403 148 407
rect 162 403 164 411
rect 118 398 120 401
rect 128 398 130 402
rect 138 401 148 403
rect 154 401 167 403
rect 138 398 140 401
rect 154 398 156 401
rect 165 400 167 401
rect 182 400 184 413
rect 189 408 191 413
rect 202 408 204 413
rect 281 425 283 433
rect 291 425 293 429
rect 304 425 306 433
rect 304 423 309 425
rect 327 424 329 429
rect 334 424 336 429
rect 307 420 309 423
rect 188 406 194 408
rect 188 404 190 406
rect 192 404 194 406
rect 188 402 194 404
rect 198 406 204 408
rect 198 404 200 406
rect 202 404 204 406
rect 198 402 204 404
rect 165 398 171 400
rect 78 373 80 378
rect 88 373 90 378
rect 98 376 100 380
rect 50 367 52 371
rect 128 376 130 380
rect 138 376 140 380
rect 118 367 120 371
rect 165 396 167 398
rect 169 396 171 398
rect 165 394 171 396
rect 178 398 184 400
rect 178 396 180 398
rect 182 396 184 398
rect 178 394 184 396
rect 182 391 184 394
rect 192 391 194 402
rect 202 398 204 402
rect 222 401 224 411
rect 232 408 234 411
rect 242 408 244 411
rect 228 406 234 408
rect 228 404 230 406
rect 232 404 234 406
rect 228 402 234 404
rect 238 406 244 408
rect 264 407 266 416
rect 271 413 273 416
rect 271 411 275 413
rect 281 412 283 416
rect 291 413 293 416
rect 273 408 275 411
rect 291 411 300 413
rect 347 422 349 426
rect 410 433 435 435
rect 410 425 412 433
rect 423 425 425 429
rect 433 425 435 433
rect 443 428 445 433
rect 450 428 452 433
rect 367 417 369 422
rect 377 417 379 422
rect 387 420 389 425
rect 407 423 412 425
rect 407 420 409 423
rect 291 409 296 411
rect 298 409 300 411
rect 238 404 240 406
rect 242 404 244 406
rect 238 402 244 404
rect 218 399 224 401
rect 218 397 220 399
rect 222 397 224 399
rect 218 395 224 397
rect 222 392 224 395
rect 229 392 231 402
rect 242 399 244 402
rect 263 405 269 407
rect 263 403 265 405
rect 267 403 269 405
rect 263 401 269 403
rect 273 406 279 408
rect 273 404 275 406
rect 277 404 279 406
rect 273 402 279 404
rect 291 407 300 409
rect 291 403 293 407
rect 307 403 309 411
rect 182 373 184 378
rect 192 373 194 378
rect 202 376 204 380
rect 154 367 156 371
rect 263 398 265 401
rect 273 398 275 402
rect 283 401 293 403
rect 299 401 312 403
rect 283 398 285 401
rect 299 398 301 401
rect 310 400 312 401
rect 327 400 329 413
rect 334 408 336 413
rect 347 408 349 413
rect 471 433 490 435
rect 471 423 473 433
rect 481 425 483 429
rect 488 425 490 433
rect 535 433 554 435
rect 498 425 500 430
rect 505 425 507 430
rect 515 425 517 430
rect 423 413 425 416
rect 416 411 425 413
rect 433 412 435 416
rect 443 413 445 416
rect 333 406 339 408
rect 333 404 335 406
rect 337 404 339 406
rect 333 402 339 404
rect 343 406 349 408
rect 343 404 345 406
rect 347 404 349 406
rect 343 402 349 404
rect 310 398 316 400
rect 242 376 244 381
rect 222 367 224 371
rect 229 367 231 371
rect 273 376 275 380
rect 283 376 285 380
rect 263 367 265 371
rect 310 396 312 398
rect 314 396 316 398
rect 310 394 316 396
rect 323 398 329 400
rect 323 396 325 398
rect 327 396 329 398
rect 323 394 329 396
rect 327 391 329 394
rect 337 391 339 402
rect 347 398 349 402
rect 367 401 369 411
rect 377 408 379 411
rect 387 408 389 411
rect 373 406 379 408
rect 373 404 375 406
rect 377 404 379 406
rect 373 402 379 404
rect 383 406 389 408
rect 383 404 385 406
rect 387 404 389 406
rect 383 402 389 404
rect 407 403 409 411
rect 416 409 418 411
rect 420 409 425 411
rect 416 407 425 409
rect 441 411 445 413
rect 441 408 443 411
rect 423 403 425 407
rect 437 406 443 408
rect 450 407 452 416
rect 437 404 439 406
rect 441 404 443 406
rect 363 399 369 401
rect 363 397 365 399
rect 367 397 369 399
rect 363 395 369 397
rect 367 392 369 395
rect 374 392 376 402
rect 387 399 389 402
rect 404 401 417 403
rect 423 401 433 403
rect 437 402 443 404
rect 404 400 406 401
rect 327 373 329 378
rect 337 373 339 378
rect 347 376 349 380
rect 299 367 301 371
rect 400 398 406 400
rect 415 398 417 401
rect 431 398 433 401
rect 441 398 443 402
rect 447 405 453 407
rect 447 403 449 405
rect 451 403 453 405
rect 447 401 453 403
rect 451 398 453 401
rect 471 399 473 417
rect 481 408 483 417
rect 477 406 483 408
rect 477 404 479 406
rect 481 404 483 406
rect 477 402 483 404
rect 488 404 490 417
rect 498 414 500 417
rect 494 412 500 414
rect 494 410 496 412
rect 498 410 500 412
rect 494 408 500 410
rect 488 402 500 404
rect 505 403 507 417
rect 535 423 537 433
rect 545 425 547 429
rect 552 425 554 433
rect 599 433 618 435
rect 562 425 564 430
rect 569 425 571 430
rect 579 425 581 430
rect 515 413 517 416
rect 512 411 518 413
rect 512 409 514 411
rect 516 409 518 411
rect 512 407 518 409
rect 400 396 402 398
rect 404 396 406 398
rect 400 394 406 396
rect 387 376 389 381
rect 367 367 369 371
rect 374 367 376 371
rect 431 376 433 380
rect 441 376 443 380
rect 415 367 417 371
rect 471 388 473 391
rect 464 386 473 388
rect 481 387 483 402
rect 487 396 493 398
rect 487 394 489 396
rect 491 394 493 396
rect 487 392 493 394
rect 488 387 490 392
rect 498 387 500 402
rect 504 401 510 403
rect 504 399 506 401
rect 508 399 510 401
rect 504 397 510 399
rect 505 387 507 397
rect 515 389 517 407
rect 535 399 537 417
rect 545 408 547 417
rect 541 406 547 408
rect 541 404 543 406
rect 545 404 547 406
rect 541 402 547 404
rect 552 404 554 417
rect 562 414 564 417
rect 558 412 564 414
rect 558 410 560 412
rect 562 410 564 412
rect 558 408 564 410
rect 552 402 564 404
rect 569 403 571 417
rect 599 423 601 433
rect 609 425 611 429
rect 616 425 618 433
rect 626 425 628 430
rect 633 425 635 430
rect 643 425 645 430
rect 579 413 581 416
rect 576 411 582 413
rect 576 409 578 411
rect 580 409 582 411
rect 576 407 582 409
rect 464 384 466 386
rect 468 384 470 386
rect 464 382 470 384
rect 535 388 537 391
rect 528 386 537 388
rect 545 387 547 402
rect 551 396 557 398
rect 551 394 553 396
rect 555 394 557 396
rect 551 392 557 394
rect 552 387 554 392
rect 562 387 564 402
rect 568 401 574 403
rect 568 399 570 401
rect 572 399 574 401
rect 568 397 574 399
rect 569 387 571 397
rect 579 389 581 407
rect 599 399 601 417
rect 609 408 611 417
rect 605 406 611 408
rect 605 404 607 406
rect 609 404 611 406
rect 605 402 611 404
rect 616 404 618 417
rect 626 414 628 417
rect 622 412 628 414
rect 622 410 624 412
rect 626 410 628 412
rect 622 408 628 410
rect 616 402 628 404
rect 633 403 635 417
rect 643 413 645 416
rect 640 411 646 413
rect 640 409 642 411
rect 644 409 646 411
rect 640 407 646 409
rect 528 384 530 386
rect 532 384 534 386
rect 528 382 534 384
rect 599 388 601 391
rect 592 386 601 388
rect 609 387 611 402
rect 615 396 621 398
rect 615 394 617 396
rect 619 394 621 396
rect 615 392 621 394
rect 616 387 618 392
rect 626 387 628 402
rect 632 401 638 403
rect 632 399 634 401
rect 636 399 638 401
rect 632 397 638 399
rect 633 387 635 397
rect 643 389 645 407
rect 592 384 594 386
rect 596 384 598 386
rect 592 382 598 384
rect 451 367 453 371
rect 481 367 483 371
rect 488 367 490 371
rect 498 367 500 371
rect 505 367 507 371
rect 515 367 517 371
rect 545 367 547 371
rect 552 367 554 371
rect 562 367 564 371
rect 569 367 571 371
rect 579 367 581 371
rect 609 367 611 371
rect 616 367 618 371
rect 626 367 628 371
rect 633 367 635 371
rect 643 367 645 371
rect 27 359 29 363
rect 34 359 36 363
rect 14 349 16 354
rect 102 359 104 363
rect 54 350 56 354
rect 64 352 66 357
rect 74 352 76 357
rect 14 328 16 331
rect 27 328 29 338
rect 34 335 36 338
rect 34 333 40 335
rect 34 331 36 333
rect 38 331 40 333
rect 34 329 40 331
rect 14 326 20 328
rect 14 324 16 326
rect 18 324 20 326
rect 14 322 20 324
rect 24 326 30 328
rect 24 324 26 326
rect 28 324 30 326
rect 24 322 30 324
rect 14 319 16 322
rect 24 319 26 322
rect 34 319 36 329
rect 54 328 56 332
rect 64 328 66 339
rect 74 336 76 339
rect 74 334 80 336
rect 74 332 76 334
rect 78 332 80 334
rect 74 330 80 332
rect 87 334 93 336
rect 87 332 89 334
rect 91 332 93 334
rect 138 359 140 363
rect 118 350 120 354
rect 128 350 130 354
rect 206 359 208 363
rect 158 350 160 354
rect 168 352 170 357
rect 178 352 180 357
rect 87 330 93 332
rect 54 326 60 328
rect 54 324 56 326
rect 58 324 60 326
rect 54 322 60 324
rect 64 326 70 328
rect 64 324 66 326
rect 68 324 70 326
rect 64 322 70 324
rect 54 317 56 322
rect 67 317 69 322
rect 74 317 76 330
rect 91 329 93 330
rect 102 329 104 332
rect 118 329 120 332
rect 91 327 104 329
rect 110 327 120 329
rect 128 328 130 332
rect 138 329 140 332
rect 94 319 96 327
rect 110 323 112 327
rect 103 321 112 323
rect 124 326 130 328
rect 124 324 126 326
rect 128 324 130 326
rect 124 322 130 324
rect 134 327 140 329
rect 134 325 136 327
rect 138 325 140 327
rect 134 323 140 325
rect 158 328 160 332
rect 168 328 170 339
rect 178 336 180 339
rect 178 334 184 336
rect 178 332 180 334
rect 182 332 184 334
rect 178 330 184 332
rect 191 334 197 336
rect 191 332 193 334
rect 195 332 197 334
rect 242 359 244 363
rect 263 359 265 363
rect 222 350 224 354
rect 232 350 234 354
rect 299 359 301 363
rect 273 350 275 354
rect 283 350 285 354
rect 367 359 369 363
rect 374 359 376 363
rect 327 352 329 357
rect 337 352 339 357
rect 347 350 349 354
rect 327 336 329 339
rect 310 334 316 336
rect 310 332 312 334
rect 314 332 316 334
rect 191 330 197 332
rect 158 326 164 328
rect 158 324 160 326
rect 162 324 164 326
rect 103 319 105 321
rect 107 319 112 321
rect 14 305 16 310
rect 24 308 26 313
rect 34 308 36 313
rect 54 304 56 308
rect 103 317 112 319
rect 128 319 130 322
rect 110 314 112 317
rect 120 314 122 318
rect 128 317 132 319
rect 130 314 132 317
rect 137 314 139 323
rect 158 322 164 324
rect 168 326 174 328
rect 168 324 170 326
rect 172 324 174 326
rect 168 322 174 324
rect 158 317 160 322
rect 171 317 173 322
rect 178 317 180 330
rect 195 329 197 330
rect 206 329 208 332
rect 222 329 224 332
rect 195 327 208 329
rect 214 327 224 329
rect 232 328 234 332
rect 242 329 244 332
rect 198 319 200 327
rect 214 323 216 327
rect 207 321 216 323
rect 228 326 234 328
rect 228 324 230 326
rect 232 324 234 326
rect 228 322 234 324
rect 238 327 244 329
rect 238 325 240 327
rect 242 325 244 327
rect 238 323 244 325
rect 263 329 265 332
rect 263 327 269 329
rect 263 325 265 327
rect 267 325 269 327
rect 263 323 269 325
rect 273 328 275 332
rect 283 329 285 332
rect 299 329 301 332
rect 310 330 316 332
rect 323 334 329 336
rect 323 332 325 334
rect 327 332 329 334
rect 323 330 329 332
rect 310 329 312 330
rect 273 326 279 328
rect 283 327 293 329
rect 299 327 312 329
rect 273 324 275 326
rect 277 324 279 326
rect 207 319 209 321
rect 211 319 216 321
rect 94 307 96 310
rect 67 301 69 306
rect 74 301 76 306
rect 94 305 99 307
rect 97 297 99 305
rect 110 301 112 305
rect 120 297 122 305
rect 158 304 160 308
rect 207 317 216 319
rect 232 319 234 322
rect 214 314 216 317
rect 224 314 226 318
rect 232 317 236 319
rect 234 314 236 317
rect 241 314 243 323
rect 264 314 266 323
rect 273 322 279 324
rect 291 323 293 327
rect 273 319 275 322
rect 271 317 275 319
rect 291 321 300 323
rect 291 319 296 321
rect 298 319 300 321
rect 307 319 309 327
rect 271 314 273 317
rect 281 314 283 318
rect 291 317 300 319
rect 291 314 293 317
rect 198 307 200 310
rect 130 297 132 302
rect 137 297 139 302
rect 97 295 122 297
rect 171 301 173 306
rect 178 301 180 306
rect 198 305 203 307
rect 201 297 203 305
rect 214 301 216 305
rect 224 297 226 305
rect 234 297 236 302
rect 241 297 243 302
rect 201 295 226 297
rect 327 317 329 330
rect 337 328 339 339
rect 415 359 417 363
rect 387 349 389 354
rect 367 335 369 338
rect 363 333 369 335
rect 347 328 349 332
rect 363 331 365 333
rect 367 331 369 333
rect 363 329 369 331
rect 333 326 339 328
rect 333 324 335 326
rect 337 324 339 326
rect 333 322 339 324
rect 343 326 349 328
rect 343 324 345 326
rect 347 324 349 326
rect 343 322 349 324
rect 334 317 336 322
rect 347 317 349 322
rect 367 319 369 329
rect 374 328 376 338
rect 400 334 406 336
rect 400 332 402 334
rect 404 332 406 334
rect 451 359 453 363
rect 481 359 483 363
rect 488 359 490 363
rect 498 359 500 363
rect 505 359 507 363
rect 515 359 517 363
rect 545 359 547 363
rect 552 359 554 363
rect 562 359 564 363
rect 569 359 571 363
rect 579 359 581 363
rect 609 359 611 363
rect 616 359 618 363
rect 626 359 628 363
rect 633 359 635 363
rect 643 359 645 363
rect 431 350 433 354
rect 441 350 443 354
rect 464 346 470 348
rect 464 344 466 346
rect 468 344 470 346
rect 464 342 473 344
rect 471 339 473 342
rect 387 328 389 331
rect 400 330 406 332
rect 373 326 379 328
rect 373 324 375 326
rect 377 324 379 326
rect 373 322 379 324
rect 383 326 389 328
rect 404 329 406 330
rect 415 329 417 332
rect 431 329 433 332
rect 404 327 417 329
rect 423 327 433 329
rect 441 328 443 332
rect 451 329 453 332
rect 383 324 385 326
rect 387 324 389 326
rect 383 322 389 324
rect 377 319 379 322
rect 387 319 389 322
rect 407 319 409 327
rect 423 323 425 327
rect 416 321 425 323
rect 437 326 443 328
rect 437 324 439 326
rect 441 324 443 326
rect 437 322 443 324
rect 447 327 453 329
rect 447 325 449 327
rect 451 325 453 327
rect 447 323 453 325
rect 416 319 418 321
rect 420 319 425 321
rect 307 307 309 310
rect 304 305 309 307
rect 264 297 266 302
rect 271 297 273 302
rect 281 297 283 305
rect 291 301 293 305
rect 304 297 306 305
rect 281 295 306 297
rect 327 301 329 306
rect 334 301 336 306
rect 347 304 349 308
rect 367 308 369 313
rect 377 308 379 313
rect 416 317 425 319
rect 441 319 443 322
rect 423 314 425 317
rect 433 314 435 318
rect 441 317 445 319
rect 443 314 445 317
rect 450 314 452 323
rect 387 305 389 310
rect 407 307 409 310
rect 407 305 412 307
rect 410 297 412 305
rect 423 301 425 305
rect 433 297 435 305
rect 471 313 473 331
rect 481 328 483 343
rect 488 338 490 343
rect 487 336 493 338
rect 487 334 489 336
rect 491 334 493 336
rect 487 332 493 334
rect 498 328 500 343
rect 505 333 507 343
rect 528 346 534 348
rect 528 344 530 346
rect 532 344 534 346
rect 528 342 537 344
rect 477 326 483 328
rect 477 324 479 326
rect 481 324 483 326
rect 477 322 483 324
rect 481 313 483 322
rect 488 326 500 328
rect 504 331 510 333
rect 504 329 506 331
rect 508 329 510 331
rect 504 327 510 329
rect 488 313 490 326
rect 494 320 500 322
rect 494 318 496 320
rect 498 318 500 320
rect 494 316 500 318
rect 498 313 500 316
rect 505 313 507 327
rect 515 323 517 341
rect 535 339 537 342
rect 512 321 518 323
rect 512 319 514 321
rect 516 319 518 321
rect 512 317 518 319
rect 515 314 517 317
rect 443 297 445 302
rect 450 297 452 302
rect 410 295 435 297
rect 471 297 473 307
rect 535 313 537 331
rect 545 328 547 343
rect 552 338 554 343
rect 551 336 557 338
rect 551 334 553 336
rect 555 334 557 336
rect 551 332 557 334
rect 562 328 564 343
rect 569 333 571 343
rect 592 346 598 348
rect 592 344 594 346
rect 596 344 598 346
rect 592 342 601 344
rect 541 326 547 328
rect 541 324 543 326
rect 545 324 547 326
rect 541 322 547 324
rect 545 313 547 322
rect 552 326 564 328
rect 568 331 574 333
rect 568 329 570 331
rect 572 329 574 331
rect 568 327 574 329
rect 552 313 554 326
rect 558 320 564 322
rect 558 318 560 320
rect 562 318 564 320
rect 558 316 564 318
rect 562 313 564 316
rect 569 313 571 327
rect 579 323 581 341
rect 599 339 601 342
rect 576 321 582 323
rect 576 319 578 321
rect 580 319 582 321
rect 576 317 582 319
rect 579 314 581 317
rect 481 301 483 305
rect 488 297 490 305
rect 498 300 500 305
rect 505 300 507 305
rect 515 300 517 305
rect 471 295 490 297
rect 535 297 537 307
rect 599 313 601 331
rect 609 328 611 343
rect 616 338 618 343
rect 615 336 621 338
rect 615 334 617 336
rect 619 334 621 336
rect 615 332 621 334
rect 626 328 628 343
rect 633 333 635 343
rect 605 326 611 328
rect 605 324 607 326
rect 609 324 611 326
rect 605 322 611 324
rect 609 313 611 322
rect 616 326 628 328
rect 632 331 638 333
rect 632 329 634 331
rect 636 329 638 331
rect 632 327 638 329
rect 616 313 618 326
rect 622 320 628 322
rect 622 318 624 320
rect 626 318 628 320
rect 622 316 628 318
rect 626 313 628 316
rect 633 313 635 327
rect 643 323 645 341
rect 640 321 646 323
rect 640 319 642 321
rect 644 319 646 321
rect 640 317 646 319
rect 643 314 645 317
rect 545 301 547 305
rect 552 297 554 305
rect 562 300 564 305
rect 569 300 571 305
rect 579 300 581 305
rect 535 295 554 297
rect 599 297 601 307
rect 609 301 611 305
rect 616 297 618 305
rect 626 300 628 305
rect 633 300 635 305
rect 643 300 645 305
rect 599 295 618 297
rect 32 289 57 291
rect 15 284 17 289
rect 22 284 24 289
rect 32 281 34 289
rect 42 281 44 285
rect 55 281 57 289
rect 55 279 60 281
rect 78 280 80 285
rect 85 280 87 285
rect 136 289 161 291
rect 119 284 121 289
rect 126 284 128 289
rect 58 276 60 279
rect 15 263 17 272
rect 22 269 24 272
rect 22 267 26 269
rect 32 268 34 272
rect 42 269 44 272
rect 24 264 26 267
rect 42 267 51 269
rect 98 278 100 282
rect 136 281 138 289
rect 146 281 148 285
rect 159 281 161 289
rect 159 279 164 281
rect 182 280 184 285
rect 189 280 191 285
rect 162 276 164 279
rect 42 265 47 267
rect 49 265 51 267
rect 14 261 20 263
rect 14 259 16 261
rect 18 259 20 261
rect 14 257 20 259
rect 24 262 30 264
rect 24 260 26 262
rect 28 260 30 262
rect 24 258 30 260
rect 42 263 51 265
rect 42 259 44 263
rect 58 259 60 267
rect 14 254 16 257
rect 24 254 26 258
rect 34 257 44 259
rect 50 257 63 259
rect 34 254 36 257
rect 50 254 52 257
rect 61 256 63 257
rect 78 256 80 269
rect 85 264 87 269
rect 98 264 100 269
rect 84 262 90 264
rect 84 260 86 262
rect 88 260 90 262
rect 84 258 90 260
rect 94 262 100 264
rect 119 263 121 272
rect 126 269 128 272
rect 126 267 130 269
rect 136 268 138 272
rect 146 269 148 272
rect 128 264 130 267
rect 146 267 155 269
rect 202 278 204 282
rect 281 289 306 291
rect 264 284 266 289
rect 271 284 273 289
rect 222 273 224 278
rect 232 273 234 278
rect 242 276 244 281
rect 146 265 151 267
rect 153 265 155 267
rect 94 260 96 262
rect 98 260 100 262
rect 94 258 100 260
rect 61 254 67 256
rect 24 232 26 236
rect 34 232 36 236
rect 14 223 16 227
rect 61 252 63 254
rect 65 252 67 254
rect 61 250 67 252
rect 74 254 80 256
rect 74 252 76 254
rect 78 252 80 254
rect 74 250 80 252
rect 78 247 80 250
rect 88 247 90 258
rect 98 254 100 258
rect 118 261 124 263
rect 118 259 120 261
rect 122 259 124 261
rect 118 257 124 259
rect 128 262 134 264
rect 128 260 130 262
rect 132 260 134 262
rect 128 258 134 260
rect 146 263 155 265
rect 146 259 148 263
rect 162 259 164 267
rect 118 254 120 257
rect 128 254 130 258
rect 138 257 148 259
rect 154 257 167 259
rect 138 254 140 257
rect 154 254 156 257
rect 165 256 167 257
rect 182 256 184 269
rect 189 264 191 269
rect 202 264 204 269
rect 281 281 283 289
rect 291 281 293 285
rect 304 281 306 289
rect 304 279 309 281
rect 327 280 329 285
rect 334 280 336 285
rect 307 276 309 279
rect 188 262 194 264
rect 188 260 190 262
rect 192 260 194 262
rect 188 258 194 260
rect 198 262 204 264
rect 198 260 200 262
rect 202 260 204 262
rect 198 258 204 260
rect 165 254 171 256
rect 78 229 80 234
rect 88 229 90 234
rect 98 232 100 236
rect 50 223 52 227
rect 128 232 130 236
rect 138 232 140 236
rect 118 223 120 227
rect 165 252 167 254
rect 169 252 171 254
rect 165 250 171 252
rect 178 254 184 256
rect 178 252 180 254
rect 182 252 184 254
rect 178 250 184 252
rect 182 247 184 250
rect 192 247 194 258
rect 202 254 204 258
rect 222 257 224 267
rect 232 264 234 267
rect 242 264 244 267
rect 228 262 234 264
rect 228 260 230 262
rect 232 260 234 262
rect 228 258 234 260
rect 238 262 244 264
rect 264 263 266 272
rect 271 269 273 272
rect 271 267 275 269
rect 281 268 283 272
rect 291 269 293 272
rect 273 264 275 267
rect 291 267 300 269
rect 347 278 349 282
rect 410 289 435 291
rect 410 281 412 289
rect 423 281 425 285
rect 433 281 435 289
rect 443 284 445 289
rect 450 284 452 289
rect 367 273 369 278
rect 377 273 379 278
rect 387 276 389 281
rect 407 279 412 281
rect 407 276 409 279
rect 291 265 296 267
rect 298 265 300 267
rect 238 260 240 262
rect 242 260 244 262
rect 238 258 244 260
rect 218 255 224 257
rect 218 253 220 255
rect 222 253 224 255
rect 218 251 224 253
rect 222 248 224 251
rect 229 248 231 258
rect 242 255 244 258
rect 263 261 269 263
rect 263 259 265 261
rect 267 259 269 261
rect 263 257 269 259
rect 273 262 279 264
rect 273 260 275 262
rect 277 260 279 262
rect 273 258 279 260
rect 291 263 300 265
rect 291 259 293 263
rect 307 259 309 267
rect 182 229 184 234
rect 192 229 194 234
rect 202 232 204 236
rect 154 223 156 227
rect 263 254 265 257
rect 273 254 275 258
rect 283 257 293 259
rect 299 257 312 259
rect 283 254 285 257
rect 299 254 301 257
rect 310 256 312 257
rect 327 256 329 269
rect 334 264 336 269
rect 347 264 349 269
rect 471 289 490 291
rect 471 279 473 289
rect 481 281 483 285
rect 488 281 490 289
rect 535 289 554 291
rect 498 281 500 286
rect 505 281 507 286
rect 515 281 517 286
rect 423 269 425 272
rect 416 267 425 269
rect 433 268 435 272
rect 443 269 445 272
rect 333 262 339 264
rect 333 260 335 262
rect 337 260 339 262
rect 333 258 339 260
rect 343 262 349 264
rect 343 260 345 262
rect 347 260 349 262
rect 343 258 349 260
rect 310 254 316 256
rect 242 232 244 237
rect 222 223 224 227
rect 229 223 231 227
rect 273 232 275 236
rect 283 232 285 236
rect 263 223 265 227
rect 310 252 312 254
rect 314 252 316 254
rect 310 250 316 252
rect 323 254 329 256
rect 323 252 325 254
rect 327 252 329 254
rect 323 250 329 252
rect 327 247 329 250
rect 337 247 339 258
rect 347 254 349 258
rect 367 257 369 267
rect 377 264 379 267
rect 387 264 389 267
rect 373 262 379 264
rect 373 260 375 262
rect 377 260 379 262
rect 373 258 379 260
rect 383 262 389 264
rect 383 260 385 262
rect 387 260 389 262
rect 383 258 389 260
rect 407 259 409 267
rect 416 265 418 267
rect 420 265 425 267
rect 416 263 425 265
rect 441 267 445 269
rect 441 264 443 267
rect 423 259 425 263
rect 437 262 443 264
rect 450 263 452 272
rect 437 260 439 262
rect 441 260 443 262
rect 363 255 369 257
rect 363 253 365 255
rect 367 253 369 255
rect 363 251 369 253
rect 367 248 369 251
rect 374 248 376 258
rect 387 255 389 258
rect 404 257 417 259
rect 423 257 433 259
rect 437 258 443 260
rect 404 256 406 257
rect 327 229 329 234
rect 337 229 339 234
rect 347 232 349 236
rect 299 223 301 227
rect 400 254 406 256
rect 415 254 417 257
rect 431 254 433 257
rect 441 254 443 258
rect 447 261 453 263
rect 447 259 449 261
rect 451 259 453 261
rect 447 257 453 259
rect 451 254 453 257
rect 471 255 473 273
rect 481 264 483 273
rect 477 262 483 264
rect 477 260 479 262
rect 481 260 483 262
rect 477 258 483 260
rect 488 260 490 273
rect 498 270 500 273
rect 494 268 500 270
rect 494 266 496 268
rect 498 266 500 268
rect 494 264 500 266
rect 488 258 500 260
rect 505 259 507 273
rect 535 279 537 289
rect 545 281 547 285
rect 552 281 554 289
rect 599 289 618 291
rect 562 281 564 286
rect 569 281 571 286
rect 579 281 581 286
rect 515 269 517 272
rect 512 267 518 269
rect 512 265 514 267
rect 516 265 518 267
rect 512 263 518 265
rect 400 252 402 254
rect 404 252 406 254
rect 400 250 406 252
rect 387 232 389 237
rect 367 223 369 227
rect 374 223 376 227
rect 431 232 433 236
rect 441 232 443 236
rect 415 223 417 227
rect 471 244 473 247
rect 464 242 473 244
rect 481 243 483 258
rect 487 252 493 254
rect 487 250 489 252
rect 491 250 493 252
rect 487 248 493 250
rect 488 243 490 248
rect 498 243 500 258
rect 504 257 510 259
rect 504 255 506 257
rect 508 255 510 257
rect 504 253 510 255
rect 505 243 507 253
rect 515 245 517 263
rect 535 255 537 273
rect 545 264 547 273
rect 541 262 547 264
rect 541 260 543 262
rect 545 260 547 262
rect 541 258 547 260
rect 552 260 554 273
rect 562 270 564 273
rect 558 268 564 270
rect 558 266 560 268
rect 562 266 564 268
rect 558 264 564 266
rect 552 258 564 260
rect 569 259 571 273
rect 599 279 601 289
rect 609 281 611 285
rect 616 281 618 289
rect 626 281 628 286
rect 633 281 635 286
rect 643 281 645 286
rect 579 269 581 272
rect 576 267 582 269
rect 576 265 578 267
rect 580 265 582 267
rect 576 263 582 265
rect 464 240 466 242
rect 468 240 470 242
rect 464 238 470 240
rect 535 244 537 247
rect 528 242 537 244
rect 545 243 547 258
rect 551 252 557 254
rect 551 250 553 252
rect 555 250 557 252
rect 551 248 557 250
rect 552 243 554 248
rect 562 243 564 258
rect 568 257 574 259
rect 568 255 570 257
rect 572 255 574 257
rect 568 253 574 255
rect 569 243 571 253
rect 579 245 581 263
rect 599 255 601 273
rect 609 264 611 273
rect 605 262 611 264
rect 605 260 607 262
rect 609 260 611 262
rect 605 258 611 260
rect 616 260 618 273
rect 626 270 628 273
rect 622 268 628 270
rect 622 266 624 268
rect 626 266 628 268
rect 622 264 628 266
rect 616 258 628 260
rect 633 259 635 273
rect 643 269 645 272
rect 640 267 646 269
rect 640 265 642 267
rect 644 265 646 267
rect 640 263 646 265
rect 528 240 530 242
rect 532 240 534 242
rect 528 238 534 240
rect 599 244 601 247
rect 592 242 601 244
rect 609 243 611 258
rect 615 252 621 254
rect 615 250 617 252
rect 619 250 621 252
rect 615 248 621 250
rect 616 243 618 248
rect 626 243 628 258
rect 632 257 638 259
rect 632 255 634 257
rect 636 255 638 257
rect 632 253 638 255
rect 633 243 635 253
rect 643 245 645 263
rect 592 240 594 242
rect 596 240 598 242
rect 592 238 598 240
rect 451 223 453 227
rect 481 223 483 227
rect 488 223 490 227
rect 498 223 500 227
rect 505 223 507 227
rect 515 223 517 227
rect 545 223 547 227
rect 552 223 554 227
rect 562 223 564 227
rect 569 223 571 227
rect 579 223 581 227
rect 609 223 611 227
rect 616 223 618 227
rect 626 223 628 227
rect 633 223 635 227
rect 643 223 645 227
rect 27 215 29 219
rect 34 215 36 219
rect 14 205 16 210
rect 102 215 104 219
rect 54 206 56 210
rect 64 208 66 213
rect 74 208 76 213
rect 14 184 16 187
rect 27 184 29 194
rect 34 191 36 194
rect 34 189 40 191
rect 34 187 36 189
rect 38 187 40 189
rect 34 185 40 187
rect 14 182 20 184
rect 14 180 16 182
rect 18 180 20 182
rect 14 178 20 180
rect 24 182 30 184
rect 24 180 26 182
rect 28 180 30 182
rect 24 178 30 180
rect 14 175 16 178
rect 24 175 26 178
rect 34 175 36 185
rect 54 184 56 188
rect 64 184 66 195
rect 74 192 76 195
rect 74 190 80 192
rect 74 188 76 190
rect 78 188 80 190
rect 74 186 80 188
rect 87 190 93 192
rect 87 188 89 190
rect 91 188 93 190
rect 138 215 140 219
rect 118 206 120 210
rect 128 206 130 210
rect 206 215 208 219
rect 158 206 160 210
rect 168 208 170 213
rect 178 208 180 213
rect 87 186 93 188
rect 54 182 60 184
rect 54 180 56 182
rect 58 180 60 182
rect 54 178 60 180
rect 64 182 70 184
rect 64 180 66 182
rect 68 180 70 182
rect 64 178 70 180
rect 54 173 56 178
rect 67 173 69 178
rect 74 173 76 186
rect 91 185 93 186
rect 102 185 104 188
rect 118 185 120 188
rect 91 183 104 185
rect 110 183 120 185
rect 128 184 130 188
rect 138 185 140 188
rect 94 175 96 183
rect 110 179 112 183
rect 103 177 112 179
rect 124 182 130 184
rect 124 180 126 182
rect 128 180 130 182
rect 124 178 130 180
rect 134 183 140 185
rect 134 181 136 183
rect 138 181 140 183
rect 134 179 140 181
rect 158 184 160 188
rect 168 184 170 195
rect 178 192 180 195
rect 178 190 184 192
rect 178 188 180 190
rect 182 188 184 190
rect 178 186 184 188
rect 191 190 197 192
rect 191 188 193 190
rect 195 188 197 190
rect 242 215 244 219
rect 263 215 265 219
rect 222 206 224 210
rect 232 206 234 210
rect 299 215 301 219
rect 273 206 275 210
rect 283 206 285 210
rect 367 215 369 219
rect 374 215 376 219
rect 327 208 329 213
rect 337 208 339 213
rect 347 206 349 210
rect 327 192 329 195
rect 310 190 316 192
rect 310 188 312 190
rect 314 188 316 190
rect 191 186 197 188
rect 158 182 164 184
rect 158 180 160 182
rect 162 180 164 182
rect 103 175 105 177
rect 107 175 112 177
rect 14 161 16 166
rect 24 164 26 169
rect 34 164 36 169
rect 54 160 56 164
rect 103 173 112 175
rect 128 175 130 178
rect 110 170 112 173
rect 120 170 122 174
rect 128 173 132 175
rect 130 170 132 173
rect 137 170 139 179
rect 158 178 164 180
rect 168 182 174 184
rect 168 180 170 182
rect 172 180 174 182
rect 168 178 174 180
rect 158 173 160 178
rect 171 173 173 178
rect 178 173 180 186
rect 195 185 197 186
rect 206 185 208 188
rect 222 185 224 188
rect 195 183 208 185
rect 214 183 224 185
rect 232 184 234 188
rect 242 185 244 188
rect 198 175 200 183
rect 214 179 216 183
rect 207 177 216 179
rect 228 182 234 184
rect 228 180 230 182
rect 232 180 234 182
rect 228 178 234 180
rect 238 183 244 185
rect 238 181 240 183
rect 242 181 244 183
rect 238 179 244 181
rect 263 185 265 188
rect 263 183 269 185
rect 263 181 265 183
rect 267 181 269 183
rect 263 179 269 181
rect 273 184 275 188
rect 283 185 285 188
rect 299 185 301 188
rect 310 186 316 188
rect 323 190 329 192
rect 323 188 325 190
rect 327 188 329 190
rect 323 186 329 188
rect 310 185 312 186
rect 273 182 279 184
rect 283 183 293 185
rect 299 183 312 185
rect 273 180 275 182
rect 277 180 279 182
rect 207 175 209 177
rect 211 175 216 177
rect 94 163 96 166
rect 67 157 69 162
rect 74 157 76 162
rect 94 161 99 163
rect 97 153 99 161
rect 110 157 112 161
rect 120 153 122 161
rect 158 160 160 164
rect 207 173 216 175
rect 232 175 234 178
rect 214 170 216 173
rect 224 170 226 174
rect 232 173 236 175
rect 234 170 236 173
rect 241 170 243 179
rect 264 170 266 179
rect 273 178 279 180
rect 291 179 293 183
rect 273 175 275 178
rect 271 173 275 175
rect 291 177 300 179
rect 291 175 296 177
rect 298 175 300 177
rect 307 175 309 183
rect 271 170 273 173
rect 281 170 283 174
rect 291 173 300 175
rect 291 170 293 173
rect 198 163 200 166
rect 130 153 132 158
rect 137 153 139 158
rect 97 151 122 153
rect 171 157 173 162
rect 178 157 180 162
rect 198 161 203 163
rect 201 153 203 161
rect 214 157 216 161
rect 224 153 226 161
rect 234 153 236 158
rect 241 153 243 158
rect 201 151 226 153
rect 327 173 329 186
rect 337 184 339 195
rect 415 215 417 219
rect 387 205 389 210
rect 367 191 369 194
rect 363 189 369 191
rect 347 184 349 188
rect 363 187 365 189
rect 367 187 369 189
rect 363 185 369 187
rect 333 182 339 184
rect 333 180 335 182
rect 337 180 339 182
rect 333 178 339 180
rect 343 182 349 184
rect 343 180 345 182
rect 347 180 349 182
rect 343 178 349 180
rect 334 173 336 178
rect 347 173 349 178
rect 367 175 369 185
rect 374 184 376 194
rect 400 190 406 192
rect 400 188 402 190
rect 404 188 406 190
rect 451 215 453 219
rect 481 215 483 219
rect 488 215 490 219
rect 498 215 500 219
rect 505 215 507 219
rect 515 215 517 219
rect 545 215 547 219
rect 552 215 554 219
rect 562 215 564 219
rect 569 215 571 219
rect 579 215 581 219
rect 609 215 611 219
rect 616 215 618 219
rect 626 215 628 219
rect 633 215 635 219
rect 643 215 645 219
rect 431 206 433 210
rect 441 206 443 210
rect 464 202 470 204
rect 464 200 466 202
rect 468 200 470 202
rect 464 198 473 200
rect 471 195 473 198
rect 387 184 389 187
rect 400 186 406 188
rect 373 182 379 184
rect 373 180 375 182
rect 377 180 379 182
rect 373 178 379 180
rect 383 182 389 184
rect 404 185 406 186
rect 415 185 417 188
rect 431 185 433 188
rect 404 183 417 185
rect 423 183 433 185
rect 441 184 443 188
rect 451 185 453 188
rect 383 180 385 182
rect 387 180 389 182
rect 383 178 389 180
rect 377 175 379 178
rect 387 175 389 178
rect 407 175 409 183
rect 423 179 425 183
rect 416 177 425 179
rect 437 182 443 184
rect 437 180 439 182
rect 441 180 443 182
rect 437 178 443 180
rect 447 183 453 185
rect 447 181 449 183
rect 451 181 453 183
rect 447 179 453 181
rect 416 175 418 177
rect 420 175 425 177
rect 307 163 309 166
rect 304 161 309 163
rect 264 153 266 158
rect 271 153 273 158
rect 281 153 283 161
rect 291 157 293 161
rect 304 153 306 161
rect 281 151 306 153
rect 327 157 329 162
rect 334 157 336 162
rect 347 160 349 164
rect 367 164 369 169
rect 377 164 379 169
rect 416 173 425 175
rect 441 175 443 178
rect 423 170 425 173
rect 433 170 435 174
rect 441 173 445 175
rect 443 170 445 173
rect 450 170 452 179
rect 387 161 389 166
rect 407 163 409 166
rect 407 161 412 163
rect 410 153 412 161
rect 423 157 425 161
rect 433 153 435 161
rect 471 169 473 187
rect 481 184 483 199
rect 488 194 490 199
rect 487 192 493 194
rect 487 190 489 192
rect 491 190 493 192
rect 487 188 493 190
rect 498 184 500 199
rect 505 189 507 199
rect 528 202 534 204
rect 528 200 530 202
rect 532 200 534 202
rect 528 198 537 200
rect 477 182 483 184
rect 477 180 479 182
rect 481 180 483 182
rect 477 178 483 180
rect 481 169 483 178
rect 488 182 500 184
rect 504 187 510 189
rect 504 185 506 187
rect 508 185 510 187
rect 504 183 510 185
rect 488 169 490 182
rect 494 176 500 178
rect 494 174 496 176
rect 498 174 500 176
rect 494 172 500 174
rect 498 169 500 172
rect 505 169 507 183
rect 515 179 517 197
rect 535 195 537 198
rect 512 177 518 179
rect 512 175 514 177
rect 516 175 518 177
rect 512 173 518 175
rect 515 170 517 173
rect 443 153 445 158
rect 450 153 452 158
rect 410 151 435 153
rect 471 153 473 163
rect 535 169 537 187
rect 545 184 547 199
rect 552 194 554 199
rect 551 192 557 194
rect 551 190 553 192
rect 555 190 557 192
rect 551 188 557 190
rect 562 184 564 199
rect 569 189 571 199
rect 592 202 598 204
rect 592 200 594 202
rect 596 200 598 202
rect 592 198 601 200
rect 541 182 547 184
rect 541 180 543 182
rect 545 180 547 182
rect 541 178 547 180
rect 545 169 547 178
rect 552 182 564 184
rect 568 187 574 189
rect 568 185 570 187
rect 572 185 574 187
rect 568 183 574 185
rect 552 169 554 182
rect 558 176 564 178
rect 558 174 560 176
rect 562 174 564 176
rect 558 172 564 174
rect 562 169 564 172
rect 569 169 571 183
rect 579 179 581 197
rect 599 195 601 198
rect 576 177 582 179
rect 576 175 578 177
rect 580 175 582 177
rect 576 173 582 175
rect 579 170 581 173
rect 481 157 483 161
rect 488 153 490 161
rect 498 156 500 161
rect 505 156 507 161
rect 515 156 517 161
rect 471 151 490 153
rect 535 153 537 163
rect 599 169 601 187
rect 609 184 611 199
rect 616 194 618 199
rect 615 192 621 194
rect 615 190 617 192
rect 619 190 621 192
rect 615 188 621 190
rect 626 184 628 199
rect 633 189 635 199
rect 605 182 611 184
rect 605 180 607 182
rect 609 180 611 182
rect 605 178 611 180
rect 609 169 611 178
rect 616 182 628 184
rect 632 187 638 189
rect 632 185 634 187
rect 636 185 638 187
rect 632 183 638 185
rect 616 169 618 182
rect 622 176 628 178
rect 622 174 624 176
rect 626 174 628 176
rect 622 172 628 174
rect 626 169 628 172
rect 633 169 635 183
rect 643 179 645 197
rect 640 177 646 179
rect 640 175 642 177
rect 644 175 646 177
rect 640 173 646 175
rect 643 170 645 173
rect 545 157 547 161
rect 552 153 554 161
rect 562 156 564 161
rect 569 156 571 161
rect 579 156 581 161
rect 535 151 554 153
rect 599 153 601 163
rect 609 157 611 161
rect 616 153 618 161
rect 626 156 628 161
rect 633 156 635 161
rect 643 156 645 161
rect 599 151 618 153
rect 32 145 57 147
rect 15 140 17 145
rect 22 140 24 145
rect 32 137 34 145
rect 42 137 44 141
rect 55 137 57 145
rect 55 135 60 137
rect 78 136 80 141
rect 85 136 87 141
rect 136 145 161 147
rect 119 140 121 145
rect 126 140 128 145
rect 58 132 60 135
rect 15 119 17 128
rect 22 125 24 128
rect 22 123 26 125
rect 32 124 34 128
rect 42 125 44 128
rect 24 120 26 123
rect 42 123 51 125
rect 98 134 100 138
rect 136 137 138 145
rect 146 137 148 141
rect 159 137 161 145
rect 159 135 164 137
rect 182 136 184 141
rect 189 136 191 141
rect 162 132 164 135
rect 42 121 47 123
rect 49 121 51 123
rect 14 117 20 119
rect 14 115 16 117
rect 18 115 20 117
rect 14 113 20 115
rect 24 118 30 120
rect 24 116 26 118
rect 28 116 30 118
rect 24 114 30 116
rect 42 119 51 121
rect 42 115 44 119
rect 58 115 60 123
rect 14 110 16 113
rect 24 110 26 114
rect 34 113 44 115
rect 50 113 63 115
rect 34 110 36 113
rect 50 110 52 113
rect 61 112 63 113
rect 78 112 80 125
rect 85 120 87 125
rect 98 120 100 125
rect 84 118 90 120
rect 84 116 86 118
rect 88 116 90 118
rect 84 114 90 116
rect 94 118 100 120
rect 119 119 121 128
rect 126 125 128 128
rect 126 123 130 125
rect 136 124 138 128
rect 146 125 148 128
rect 128 120 130 123
rect 146 123 155 125
rect 202 134 204 138
rect 281 145 306 147
rect 264 140 266 145
rect 271 140 273 145
rect 222 129 224 134
rect 232 129 234 134
rect 242 132 244 137
rect 146 121 151 123
rect 153 121 155 123
rect 94 116 96 118
rect 98 116 100 118
rect 94 114 100 116
rect 61 110 67 112
rect 24 88 26 92
rect 34 88 36 92
rect 14 79 16 83
rect 61 108 63 110
rect 65 108 67 110
rect 61 106 67 108
rect 74 110 80 112
rect 74 108 76 110
rect 78 108 80 110
rect 74 106 80 108
rect 78 103 80 106
rect 88 103 90 114
rect 98 110 100 114
rect 118 117 124 119
rect 118 115 120 117
rect 122 115 124 117
rect 118 113 124 115
rect 128 118 134 120
rect 128 116 130 118
rect 132 116 134 118
rect 128 114 134 116
rect 146 119 155 121
rect 146 115 148 119
rect 162 115 164 123
rect 118 110 120 113
rect 128 110 130 114
rect 138 113 148 115
rect 154 113 167 115
rect 138 110 140 113
rect 154 110 156 113
rect 165 112 167 113
rect 182 112 184 125
rect 189 120 191 125
rect 202 120 204 125
rect 281 137 283 145
rect 291 137 293 141
rect 304 137 306 145
rect 304 135 309 137
rect 327 136 329 141
rect 334 136 336 141
rect 307 132 309 135
rect 188 118 194 120
rect 188 116 190 118
rect 192 116 194 118
rect 188 114 194 116
rect 198 118 204 120
rect 198 116 200 118
rect 202 116 204 118
rect 198 114 204 116
rect 165 110 171 112
rect 78 85 80 90
rect 88 85 90 90
rect 98 88 100 92
rect 50 79 52 83
rect 128 88 130 92
rect 138 88 140 92
rect 118 79 120 83
rect 165 108 167 110
rect 169 108 171 110
rect 165 106 171 108
rect 178 110 184 112
rect 178 108 180 110
rect 182 108 184 110
rect 178 106 184 108
rect 182 103 184 106
rect 192 103 194 114
rect 202 110 204 114
rect 222 113 224 123
rect 232 120 234 123
rect 242 120 244 123
rect 228 118 234 120
rect 228 116 230 118
rect 232 116 234 118
rect 228 114 234 116
rect 238 118 244 120
rect 264 119 266 128
rect 271 125 273 128
rect 271 123 275 125
rect 281 124 283 128
rect 291 125 293 128
rect 273 120 275 123
rect 291 123 300 125
rect 347 134 349 138
rect 410 145 435 147
rect 410 137 412 145
rect 423 137 425 141
rect 433 137 435 145
rect 443 140 445 145
rect 450 140 452 145
rect 367 129 369 134
rect 377 129 379 134
rect 387 132 389 137
rect 407 135 412 137
rect 407 132 409 135
rect 291 121 296 123
rect 298 121 300 123
rect 238 116 240 118
rect 242 116 244 118
rect 238 114 244 116
rect 218 111 224 113
rect 218 109 220 111
rect 222 109 224 111
rect 218 107 224 109
rect 222 104 224 107
rect 229 104 231 114
rect 242 111 244 114
rect 263 117 269 119
rect 263 115 265 117
rect 267 115 269 117
rect 263 113 269 115
rect 273 118 279 120
rect 273 116 275 118
rect 277 116 279 118
rect 273 114 279 116
rect 291 119 300 121
rect 291 115 293 119
rect 307 115 309 123
rect 182 85 184 90
rect 192 85 194 90
rect 202 88 204 92
rect 154 79 156 83
rect 263 110 265 113
rect 273 110 275 114
rect 283 113 293 115
rect 299 113 312 115
rect 283 110 285 113
rect 299 110 301 113
rect 310 112 312 113
rect 327 112 329 125
rect 334 120 336 125
rect 347 120 349 125
rect 471 145 490 147
rect 471 135 473 145
rect 481 137 483 141
rect 488 137 490 145
rect 535 145 554 147
rect 498 137 500 142
rect 505 137 507 142
rect 515 137 517 142
rect 423 125 425 128
rect 416 123 425 125
rect 433 124 435 128
rect 443 125 445 128
rect 333 118 339 120
rect 333 116 335 118
rect 337 116 339 118
rect 333 114 339 116
rect 343 118 349 120
rect 343 116 345 118
rect 347 116 349 118
rect 343 114 349 116
rect 310 110 316 112
rect 242 88 244 93
rect 222 79 224 83
rect 229 79 231 83
rect 273 88 275 92
rect 283 88 285 92
rect 263 79 265 83
rect 310 108 312 110
rect 314 108 316 110
rect 310 106 316 108
rect 323 110 329 112
rect 323 108 325 110
rect 327 108 329 110
rect 323 106 329 108
rect 327 103 329 106
rect 337 103 339 114
rect 347 110 349 114
rect 367 113 369 123
rect 377 120 379 123
rect 387 120 389 123
rect 373 118 379 120
rect 373 116 375 118
rect 377 116 379 118
rect 373 114 379 116
rect 383 118 389 120
rect 383 116 385 118
rect 387 116 389 118
rect 383 114 389 116
rect 407 115 409 123
rect 416 121 418 123
rect 420 121 425 123
rect 416 119 425 121
rect 441 123 445 125
rect 441 120 443 123
rect 423 115 425 119
rect 437 118 443 120
rect 450 119 452 128
rect 437 116 439 118
rect 441 116 443 118
rect 363 111 369 113
rect 363 109 365 111
rect 367 109 369 111
rect 363 107 369 109
rect 367 104 369 107
rect 374 104 376 114
rect 387 111 389 114
rect 404 113 417 115
rect 423 113 433 115
rect 437 114 443 116
rect 404 112 406 113
rect 327 85 329 90
rect 337 85 339 90
rect 347 88 349 92
rect 299 79 301 83
rect 400 110 406 112
rect 415 110 417 113
rect 431 110 433 113
rect 441 110 443 114
rect 447 117 453 119
rect 447 115 449 117
rect 451 115 453 117
rect 447 113 453 115
rect 451 110 453 113
rect 471 111 473 129
rect 481 120 483 129
rect 477 118 483 120
rect 477 116 479 118
rect 481 116 483 118
rect 477 114 483 116
rect 488 116 490 129
rect 498 126 500 129
rect 494 124 500 126
rect 494 122 496 124
rect 498 122 500 124
rect 494 120 500 122
rect 488 114 500 116
rect 505 115 507 129
rect 535 135 537 145
rect 545 137 547 141
rect 552 137 554 145
rect 599 145 618 147
rect 562 137 564 142
rect 569 137 571 142
rect 579 137 581 142
rect 515 125 517 128
rect 512 123 518 125
rect 512 121 514 123
rect 516 121 518 123
rect 512 119 518 121
rect 400 108 402 110
rect 404 108 406 110
rect 400 106 406 108
rect 387 88 389 93
rect 367 79 369 83
rect 374 79 376 83
rect 431 88 433 92
rect 441 88 443 92
rect 415 79 417 83
rect 471 100 473 103
rect 464 98 473 100
rect 481 99 483 114
rect 487 108 493 110
rect 487 106 489 108
rect 491 106 493 108
rect 487 104 493 106
rect 488 99 490 104
rect 498 99 500 114
rect 504 113 510 115
rect 504 111 506 113
rect 508 111 510 113
rect 504 109 510 111
rect 505 99 507 109
rect 515 101 517 119
rect 535 111 537 129
rect 545 120 547 129
rect 541 118 547 120
rect 541 116 543 118
rect 545 116 547 118
rect 541 114 547 116
rect 552 116 554 129
rect 562 126 564 129
rect 558 124 564 126
rect 558 122 560 124
rect 562 122 564 124
rect 558 120 564 122
rect 552 114 564 116
rect 569 115 571 129
rect 599 135 601 145
rect 609 137 611 141
rect 616 137 618 145
rect 626 137 628 142
rect 633 137 635 142
rect 643 137 645 142
rect 579 125 581 128
rect 576 123 582 125
rect 576 121 578 123
rect 580 121 582 123
rect 576 119 582 121
rect 464 96 466 98
rect 468 96 470 98
rect 464 94 470 96
rect 535 100 537 103
rect 528 98 537 100
rect 545 99 547 114
rect 551 108 557 110
rect 551 106 553 108
rect 555 106 557 108
rect 551 104 557 106
rect 552 99 554 104
rect 562 99 564 114
rect 568 113 574 115
rect 568 111 570 113
rect 572 111 574 113
rect 568 109 574 111
rect 569 99 571 109
rect 579 101 581 119
rect 599 111 601 129
rect 609 120 611 129
rect 605 118 611 120
rect 605 116 607 118
rect 609 116 611 118
rect 605 114 611 116
rect 616 116 618 129
rect 626 126 628 129
rect 622 124 628 126
rect 622 122 624 124
rect 626 122 628 124
rect 622 120 628 122
rect 616 114 628 116
rect 633 115 635 129
rect 643 125 645 128
rect 640 123 646 125
rect 640 121 642 123
rect 644 121 646 123
rect 640 119 646 121
rect 528 96 530 98
rect 532 96 534 98
rect 528 94 534 96
rect 599 100 601 103
rect 592 98 601 100
rect 609 99 611 114
rect 615 108 621 110
rect 615 106 617 108
rect 619 106 621 108
rect 615 104 621 106
rect 616 99 618 104
rect 626 99 628 114
rect 632 113 638 115
rect 632 111 634 113
rect 636 111 638 113
rect 632 109 638 111
rect 633 99 635 109
rect 643 101 645 119
rect 592 96 594 98
rect 596 96 598 98
rect 592 94 598 96
rect 451 79 453 83
rect 481 79 483 83
rect 488 79 490 83
rect 498 79 500 83
rect 505 79 507 83
rect 515 79 517 83
rect 545 79 547 83
rect 552 79 554 83
rect 562 79 564 83
rect 569 79 571 83
rect 579 79 581 83
rect 609 79 611 83
rect 616 79 618 83
rect 626 79 628 83
rect 633 79 635 83
rect 643 79 645 83
rect 27 71 29 75
rect 34 71 36 75
rect 14 61 16 66
rect 102 71 104 75
rect 54 62 56 66
rect 64 64 66 69
rect 74 64 76 69
rect 14 40 16 43
rect 27 40 29 50
rect 34 47 36 50
rect 34 45 40 47
rect 34 43 36 45
rect 38 43 40 45
rect 34 41 40 43
rect 14 38 20 40
rect 14 36 16 38
rect 18 36 20 38
rect 14 34 20 36
rect 24 38 30 40
rect 24 36 26 38
rect 28 36 30 38
rect 24 34 30 36
rect 14 31 16 34
rect 24 31 26 34
rect 34 31 36 41
rect 54 40 56 44
rect 64 40 66 51
rect 74 48 76 51
rect 74 46 80 48
rect 74 44 76 46
rect 78 44 80 46
rect 74 42 80 44
rect 87 46 93 48
rect 87 44 89 46
rect 91 44 93 46
rect 138 71 140 75
rect 118 62 120 66
rect 128 62 130 66
rect 206 71 208 75
rect 158 62 160 66
rect 168 64 170 69
rect 178 64 180 69
rect 87 42 93 44
rect 54 38 60 40
rect 54 36 56 38
rect 58 36 60 38
rect 54 34 60 36
rect 64 38 70 40
rect 64 36 66 38
rect 68 36 70 38
rect 64 34 70 36
rect 54 29 56 34
rect 67 29 69 34
rect 74 29 76 42
rect 91 41 93 42
rect 102 41 104 44
rect 118 41 120 44
rect 91 39 104 41
rect 110 39 120 41
rect 128 40 130 44
rect 138 41 140 44
rect 94 31 96 39
rect 110 35 112 39
rect 103 33 112 35
rect 124 38 130 40
rect 124 36 126 38
rect 128 36 130 38
rect 124 34 130 36
rect 134 39 140 41
rect 134 37 136 39
rect 138 37 140 39
rect 134 35 140 37
rect 158 40 160 44
rect 168 40 170 51
rect 178 48 180 51
rect 178 46 184 48
rect 178 44 180 46
rect 182 44 184 46
rect 178 42 184 44
rect 191 46 197 48
rect 191 44 193 46
rect 195 44 197 46
rect 242 71 244 75
rect 263 71 265 75
rect 222 62 224 66
rect 232 62 234 66
rect 299 71 301 75
rect 273 62 275 66
rect 283 62 285 66
rect 367 71 369 75
rect 374 71 376 75
rect 327 64 329 69
rect 337 64 339 69
rect 347 62 349 66
rect 327 48 329 51
rect 310 46 316 48
rect 310 44 312 46
rect 314 44 316 46
rect 191 42 197 44
rect 158 38 164 40
rect 158 36 160 38
rect 162 36 164 38
rect 103 31 105 33
rect 107 31 112 33
rect 14 17 16 22
rect 24 20 26 25
rect 34 20 36 25
rect 54 16 56 20
rect 103 29 112 31
rect 128 31 130 34
rect 110 26 112 29
rect 120 26 122 30
rect 128 29 132 31
rect 130 26 132 29
rect 137 26 139 35
rect 158 34 164 36
rect 168 38 174 40
rect 168 36 170 38
rect 172 36 174 38
rect 168 34 174 36
rect 158 29 160 34
rect 171 29 173 34
rect 178 29 180 42
rect 195 41 197 42
rect 206 41 208 44
rect 222 41 224 44
rect 195 39 208 41
rect 214 39 224 41
rect 232 40 234 44
rect 242 41 244 44
rect 198 31 200 39
rect 214 35 216 39
rect 207 33 216 35
rect 228 38 234 40
rect 228 36 230 38
rect 232 36 234 38
rect 228 34 234 36
rect 238 39 244 41
rect 238 37 240 39
rect 242 37 244 39
rect 238 35 244 37
rect 263 41 265 44
rect 263 39 269 41
rect 263 37 265 39
rect 267 37 269 39
rect 263 35 269 37
rect 273 40 275 44
rect 283 41 285 44
rect 299 41 301 44
rect 310 42 316 44
rect 323 46 329 48
rect 323 44 325 46
rect 327 44 329 46
rect 323 42 329 44
rect 310 41 312 42
rect 273 38 279 40
rect 283 39 293 41
rect 299 39 312 41
rect 273 36 275 38
rect 277 36 279 38
rect 207 31 209 33
rect 211 31 216 33
rect 94 19 96 22
rect 67 13 69 18
rect 74 13 76 18
rect 94 17 99 19
rect 97 9 99 17
rect 110 13 112 17
rect 120 9 122 17
rect 158 16 160 20
rect 207 29 216 31
rect 232 31 234 34
rect 214 26 216 29
rect 224 26 226 30
rect 232 29 236 31
rect 234 26 236 29
rect 241 26 243 35
rect 264 26 266 35
rect 273 34 279 36
rect 291 35 293 39
rect 273 31 275 34
rect 271 29 275 31
rect 291 33 300 35
rect 291 31 296 33
rect 298 31 300 33
rect 307 31 309 39
rect 271 26 273 29
rect 281 26 283 30
rect 291 29 300 31
rect 291 26 293 29
rect 198 19 200 22
rect 130 9 132 14
rect 137 9 139 14
rect 97 7 122 9
rect 171 13 173 18
rect 178 13 180 18
rect 198 17 203 19
rect 201 9 203 17
rect 214 13 216 17
rect 224 9 226 17
rect 234 9 236 14
rect 241 9 243 14
rect 201 7 226 9
rect 327 29 329 42
rect 337 40 339 51
rect 415 71 417 75
rect 387 61 389 66
rect 367 47 369 50
rect 363 45 369 47
rect 347 40 349 44
rect 363 43 365 45
rect 367 43 369 45
rect 363 41 369 43
rect 333 38 339 40
rect 333 36 335 38
rect 337 36 339 38
rect 333 34 339 36
rect 343 38 349 40
rect 343 36 345 38
rect 347 36 349 38
rect 343 34 349 36
rect 334 29 336 34
rect 347 29 349 34
rect 367 31 369 41
rect 374 40 376 50
rect 400 46 406 48
rect 400 44 402 46
rect 404 44 406 46
rect 451 71 453 75
rect 481 71 483 75
rect 488 71 490 75
rect 498 71 500 75
rect 505 71 507 75
rect 515 71 517 75
rect 545 71 547 75
rect 552 71 554 75
rect 562 71 564 75
rect 569 71 571 75
rect 579 71 581 75
rect 609 71 611 75
rect 616 71 618 75
rect 626 71 628 75
rect 633 71 635 75
rect 643 71 645 75
rect 431 62 433 66
rect 441 62 443 66
rect 464 58 470 60
rect 464 56 466 58
rect 468 56 470 58
rect 464 54 473 56
rect 471 51 473 54
rect 387 40 389 43
rect 400 42 406 44
rect 373 38 379 40
rect 373 36 375 38
rect 377 36 379 38
rect 373 34 379 36
rect 383 38 389 40
rect 404 41 406 42
rect 415 41 417 44
rect 431 41 433 44
rect 404 39 417 41
rect 423 39 433 41
rect 441 40 443 44
rect 451 41 453 44
rect 383 36 385 38
rect 387 36 389 38
rect 383 34 389 36
rect 377 31 379 34
rect 387 31 389 34
rect 407 31 409 39
rect 423 35 425 39
rect 416 33 425 35
rect 437 38 443 40
rect 437 36 439 38
rect 441 36 443 38
rect 437 34 443 36
rect 447 39 453 41
rect 447 37 449 39
rect 451 37 453 39
rect 447 35 453 37
rect 416 31 418 33
rect 420 31 425 33
rect 307 19 309 22
rect 304 17 309 19
rect 264 9 266 14
rect 271 9 273 14
rect 281 9 283 17
rect 291 13 293 17
rect 304 9 306 17
rect 281 7 306 9
rect 327 13 329 18
rect 334 13 336 18
rect 347 16 349 20
rect 367 20 369 25
rect 377 20 379 25
rect 416 29 425 31
rect 441 31 443 34
rect 423 26 425 29
rect 433 26 435 30
rect 441 29 445 31
rect 443 26 445 29
rect 450 26 452 35
rect 387 17 389 22
rect 407 19 409 22
rect 407 17 412 19
rect 410 9 412 17
rect 423 13 425 17
rect 433 9 435 17
rect 471 25 473 43
rect 481 40 483 55
rect 488 50 490 55
rect 487 48 493 50
rect 487 46 489 48
rect 491 46 493 48
rect 487 44 493 46
rect 498 40 500 55
rect 505 45 507 55
rect 528 58 534 60
rect 528 56 530 58
rect 532 56 534 58
rect 528 54 537 56
rect 477 38 483 40
rect 477 36 479 38
rect 481 36 483 38
rect 477 34 483 36
rect 481 25 483 34
rect 488 38 500 40
rect 504 43 510 45
rect 504 41 506 43
rect 508 41 510 43
rect 504 39 510 41
rect 488 25 490 38
rect 494 32 500 34
rect 494 30 496 32
rect 498 30 500 32
rect 494 28 500 30
rect 498 25 500 28
rect 505 25 507 39
rect 515 35 517 53
rect 535 51 537 54
rect 512 33 518 35
rect 512 31 514 33
rect 516 31 518 33
rect 512 29 518 31
rect 515 26 517 29
rect 443 9 445 14
rect 450 9 452 14
rect 410 7 435 9
rect 471 9 473 19
rect 535 25 537 43
rect 545 40 547 55
rect 552 50 554 55
rect 551 48 557 50
rect 551 46 553 48
rect 555 46 557 48
rect 551 44 557 46
rect 562 40 564 55
rect 569 45 571 55
rect 592 58 598 60
rect 592 56 594 58
rect 596 56 598 58
rect 592 54 601 56
rect 541 38 547 40
rect 541 36 543 38
rect 545 36 547 38
rect 541 34 547 36
rect 545 25 547 34
rect 552 38 564 40
rect 568 43 574 45
rect 568 41 570 43
rect 572 41 574 43
rect 568 39 574 41
rect 552 25 554 38
rect 558 32 564 34
rect 558 30 560 32
rect 562 30 564 32
rect 558 28 564 30
rect 562 25 564 28
rect 569 25 571 39
rect 579 35 581 53
rect 599 51 601 54
rect 576 33 582 35
rect 576 31 578 33
rect 580 31 582 33
rect 576 29 582 31
rect 579 26 581 29
rect 481 13 483 17
rect 488 9 490 17
rect 498 12 500 17
rect 505 12 507 17
rect 515 12 517 17
rect 471 7 490 9
rect 535 9 537 19
rect 599 25 601 43
rect 609 40 611 55
rect 616 50 618 55
rect 615 48 621 50
rect 615 46 617 48
rect 619 46 621 48
rect 615 44 621 46
rect 626 40 628 55
rect 633 45 635 55
rect 605 38 611 40
rect 605 36 607 38
rect 609 36 611 38
rect 605 34 611 36
rect 609 25 611 34
rect 616 38 628 40
rect 632 43 638 45
rect 632 41 634 43
rect 636 41 638 43
rect 632 39 638 41
rect 616 25 618 38
rect 622 32 628 34
rect 622 30 624 32
rect 626 30 628 32
rect 622 28 628 30
rect 626 25 628 28
rect 633 25 635 39
rect 643 35 645 53
rect 640 33 646 35
rect 640 31 642 33
rect 644 31 646 33
rect 640 29 646 31
rect 643 26 645 29
rect 545 13 547 17
rect 552 9 554 17
rect 562 12 564 17
rect 569 12 571 17
rect 579 12 581 17
rect 535 7 554 9
rect 599 9 601 19
rect 609 13 611 17
rect 616 9 618 17
rect 626 12 628 17
rect 633 12 635 17
rect 643 12 645 17
rect 599 7 618 9
<< ndif >>
rect 7 576 13 578
rect 7 574 9 576
rect 11 574 13 576
rect 7 572 13 574
rect 7 560 15 572
rect 17 560 22 572
rect 24 569 29 572
rect 89 576 96 578
rect 89 574 92 576
rect 94 574 96 576
rect 24 566 32 569
rect 24 564 27 566
rect 29 564 32 566
rect 24 560 32 564
rect 34 564 42 569
rect 34 562 37 564
rect 39 562 42 564
rect 34 560 42 562
rect 44 567 53 569
rect 89 568 96 574
rect 111 576 117 578
rect 111 574 113 576
rect 115 574 117 576
rect 111 572 117 574
rect 44 565 49 567
rect 51 565 53 567
rect 44 564 53 565
rect 71 566 78 568
rect 71 564 73 566
rect 75 564 78 566
rect 44 560 58 564
rect 53 555 58 560
rect 60 561 65 564
rect 71 562 78 564
rect 60 559 67 561
rect 60 557 63 559
rect 65 557 67 559
rect 73 557 78 562
rect 80 557 85 568
rect 87 566 96 568
rect 87 557 98 566
rect 100 564 107 566
rect 100 562 103 564
rect 105 562 107 564
rect 100 560 107 562
rect 111 560 119 572
rect 121 560 126 572
rect 128 569 133 572
rect 193 576 200 578
rect 193 574 196 576
rect 198 574 200 576
rect 128 566 136 569
rect 128 564 131 566
rect 133 564 136 566
rect 128 560 136 564
rect 138 564 146 569
rect 138 562 141 564
rect 143 562 146 564
rect 138 560 146 562
rect 148 567 157 569
rect 193 568 200 574
rect 215 572 221 574
rect 215 570 217 572
rect 219 570 221 572
rect 148 565 153 567
rect 155 565 157 567
rect 148 564 157 565
rect 175 566 182 568
rect 175 564 177 566
rect 179 564 182 566
rect 148 560 162 564
rect 100 557 105 560
rect 60 555 67 557
rect 157 555 162 560
rect 164 561 169 564
rect 175 562 182 564
rect 164 559 171 561
rect 164 557 167 559
rect 169 557 171 559
rect 177 557 182 562
rect 184 557 189 568
rect 191 566 200 568
rect 215 568 221 570
rect 234 572 240 574
rect 256 576 262 578
rect 256 574 258 576
rect 260 574 262 576
rect 256 572 262 574
rect 234 570 236 572
rect 238 570 240 572
rect 234 568 240 570
rect 191 557 202 566
rect 204 564 211 566
rect 204 562 207 564
rect 209 562 211 564
rect 204 560 211 562
rect 215 561 220 568
rect 236 564 240 568
rect 236 561 242 564
rect 204 557 209 560
rect 164 555 171 557
rect 215 555 222 561
rect 224 559 232 561
rect 224 557 227 559
rect 229 557 232 559
rect 224 555 232 557
rect 234 555 242 561
rect 244 561 249 564
rect 244 559 251 561
rect 256 560 264 572
rect 266 560 271 572
rect 273 569 278 572
rect 338 576 345 578
rect 338 574 341 576
rect 343 574 345 576
rect 273 566 281 569
rect 273 564 276 566
rect 278 564 281 566
rect 273 560 281 564
rect 283 564 291 569
rect 283 562 286 564
rect 288 562 291 564
rect 283 560 291 562
rect 293 567 302 569
rect 338 568 345 574
rect 360 572 366 574
rect 360 570 362 572
rect 364 570 366 572
rect 293 565 298 567
rect 300 565 302 567
rect 293 564 302 565
rect 320 566 327 568
rect 320 564 322 566
rect 324 564 327 566
rect 293 560 307 564
rect 244 557 247 559
rect 249 557 251 559
rect 244 555 251 557
rect 302 555 307 560
rect 309 561 314 564
rect 320 562 327 564
rect 309 559 316 561
rect 309 557 312 559
rect 314 557 316 559
rect 322 557 327 562
rect 329 557 334 568
rect 336 566 345 568
rect 360 568 366 570
rect 379 572 385 574
rect 379 570 381 572
rect 383 570 385 572
rect 379 568 385 570
rect 454 576 460 578
rect 454 574 456 576
rect 458 574 460 576
rect 454 572 460 574
rect 438 569 443 572
rect 336 557 347 566
rect 349 564 356 566
rect 349 562 352 564
rect 354 562 356 564
rect 349 560 356 562
rect 360 561 365 568
rect 381 564 385 568
rect 414 567 423 569
rect 414 565 416 567
rect 418 565 423 567
rect 414 564 423 565
rect 381 561 387 564
rect 349 557 354 560
rect 309 555 316 557
rect 360 555 367 561
rect 369 559 377 561
rect 369 557 372 559
rect 374 557 377 559
rect 369 555 377 557
rect 379 555 387 561
rect 389 561 394 564
rect 402 561 407 564
rect 389 559 396 561
rect 389 557 392 559
rect 394 557 396 559
rect 389 555 396 557
rect 400 559 407 561
rect 400 557 402 559
rect 404 557 407 559
rect 400 555 407 557
rect 409 560 423 564
rect 425 564 433 569
rect 425 562 428 564
rect 430 562 433 564
rect 425 560 433 562
rect 435 566 443 569
rect 435 564 438 566
rect 440 564 443 566
rect 435 560 443 564
rect 445 560 450 572
rect 452 560 460 572
rect 475 567 481 569
rect 464 565 471 567
rect 464 563 466 565
rect 468 563 471 565
rect 464 561 471 563
rect 473 565 481 567
rect 473 563 476 565
rect 478 563 481 565
rect 473 561 481 563
rect 483 561 488 569
rect 490 567 498 569
rect 490 565 493 567
rect 495 565 498 567
rect 490 561 498 565
rect 500 561 505 569
rect 507 567 515 569
rect 507 565 510 567
rect 512 565 515 567
rect 507 561 515 565
rect 409 555 414 560
rect 510 560 515 561
rect 517 566 522 569
rect 539 567 545 569
rect 517 564 524 566
rect 517 562 520 564
rect 522 562 524 564
rect 517 560 524 562
rect 528 565 535 567
rect 528 563 530 565
rect 532 563 535 565
rect 528 561 535 563
rect 537 565 545 567
rect 537 563 540 565
rect 542 563 545 565
rect 537 561 545 563
rect 547 561 552 569
rect 554 567 562 569
rect 554 565 557 567
rect 559 565 562 567
rect 554 561 562 565
rect 564 561 569 569
rect 571 567 579 569
rect 571 565 574 567
rect 576 565 579 567
rect 571 561 579 565
rect 574 560 579 561
rect 581 566 586 569
rect 603 567 609 569
rect 581 564 588 566
rect 581 562 584 564
rect 586 562 588 564
rect 581 560 588 562
rect 592 565 599 567
rect 592 563 594 565
rect 596 563 599 565
rect 592 561 599 563
rect 601 565 609 567
rect 601 563 604 565
rect 606 563 609 565
rect 601 561 609 563
rect 611 561 616 569
rect 618 567 626 569
rect 618 565 621 567
rect 623 565 626 567
rect 618 561 626 565
rect 628 561 633 569
rect 635 567 643 569
rect 635 565 638 567
rect 640 565 643 567
rect 635 561 643 565
rect 638 560 643 561
rect 645 566 650 569
rect 645 564 652 566
rect 645 562 648 564
rect 650 562 652 564
rect 645 560 652 562
rect 7 461 14 463
rect 7 459 9 461
rect 11 459 14 461
rect 7 457 14 459
rect 9 454 14 457
rect 16 457 24 463
rect 26 461 34 463
rect 26 459 29 461
rect 31 459 34 461
rect 26 457 34 459
rect 36 457 43 463
rect 87 461 94 463
rect 49 458 54 461
rect 16 454 22 457
rect 18 450 22 454
rect 38 450 43 457
rect 47 456 54 458
rect 47 454 49 456
rect 51 454 54 456
rect 47 452 54 454
rect 56 452 67 461
rect 18 448 24 450
rect 18 446 20 448
rect 22 446 24 448
rect 18 444 24 446
rect 37 448 43 450
rect 58 450 67 452
rect 69 450 74 461
rect 76 456 81 461
rect 87 459 89 461
rect 91 459 94 461
rect 87 457 94 459
rect 76 454 83 456
rect 89 454 94 457
rect 96 458 101 463
rect 191 461 198 463
rect 153 458 158 461
rect 96 454 110 458
rect 76 452 79 454
rect 81 452 83 454
rect 76 450 83 452
rect 101 453 110 454
rect 101 451 103 453
rect 105 451 110 453
rect 37 446 39 448
rect 41 446 43 448
rect 37 444 43 446
rect 58 444 65 450
rect 101 449 110 451
rect 112 456 120 458
rect 112 454 115 456
rect 117 454 120 456
rect 112 449 120 454
rect 122 454 130 458
rect 122 452 125 454
rect 127 452 130 454
rect 122 449 130 452
rect 58 442 60 444
rect 62 442 65 444
rect 58 440 65 442
rect 125 446 130 449
rect 132 446 137 458
rect 139 446 147 458
rect 151 456 158 458
rect 151 454 153 456
rect 155 454 158 456
rect 151 452 158 454
rect 160 452 171 461
rect 162 450 171 452
rect 173 450 178 461
rect 180 456 185 461
rect 191 459 193 461
rect 195 459 198 461
rect 191 457 198 459
rect 180 454 187 456
rect 193 454 198 457
rect 200 458 205 463
rect 302 458 307 463
rect 200 454 214 458
rect 180 452 183 454
rect 185 452 187 454
rect 180 450 187 452
rect 205 453 214 454
rect 205 451 207 453
rect 209 451 214 453
rect 141 444 147 446
rect 141 442 143 444
rect 145 442 147 444
rect 141 440 147 442
rect 162 444 169 450
rect 205 449 214 451
rect 216 456 224 458
rect 216 454 219 456
rect 221 454 224 456
rect 216 449 224 454
rect 226 454 234 458
rect 226 452 229 454
rect 231 452 234 454
rect 226 449 234 452
rect 162 442 164 444
rect 166 442 169 444
rect 162 440 169 442
rect 229 446 234 449
rect 236 446 241 458
rect 243 446 251 458
rect 245 444 251 446
rect 245 442 247 444
rect 249 442 251 444
rect 245 440 251 442
rect 256 446 264 458
rect 266 446 271 458
rect 273 454 281 458
rect 273 452 276 454
rect 278 452 281 454
rect 273 449 281 452
rect 283 456 291 458
rect 283 454 286 456
rect 288 454 291 456
rect 283 449 291 454
rect 293 454 307 458
rect 309 461 316 463
rect 309 459 312 461
rect 314 459 316 461
rect 309 457 316 459
rect 309 454 314 457
rect 322 456 327 461
rect 320 454 327 456
rect 293 453 302 454
rect 293 451 298 453
rect 300 451 302 453
rect 293 449 302 451
rect 320 452 322 454
rect 324 452 327 454
rect 320 450 327 452
rect 329 450 334 461
rect 336 452 347 461
rect 349 458 354 461
rect 349 456 356 458
rect 349 454 352 456
rect 354 454 356 456
rect 349 452 356 454
rect 360 457 367 463
rect 369 461 377 463
rect 369 459 372 461
rect 374 459 377 461
rect 369 457 377 459
rect 379 457 387 463
rect 336 450 345 452
rect 273 446 278 449
rect 256 444 262 446
rect 256 442 258 444
rect 260 442 262 444
rect 256 440 262 442
rect 338 444 345 450
rect 360 450 365 457
rect 381 454 387 457
rect 389 461 396 463
rect 389 459 392 461
rect 394 459 396 461
rect 389 457 396 459
rect 400 461 407 463
rect 400 459 402 461
rect 404 459 407 461
rect 400 457 407 459
rect 389 454 394 457
rect 402 454 407 457
rect 409 458 414 463
rect 409 454 423 458
rect 381 450 385 454
rect 360 448 366 450
rect 360 446 362 448
rect 364 446 366 448
rect 338 442 341 444
rect 343 442 345 444
rect 338 440 345 442
rect 360 444 366 446
rect 379 448 385 450
rect 414 453 423 454
rect 414 451 416 453
rect 418 451 423 453
rect 414 449 423 451
rect 425 456 433 458
rect 425 454 428 456
rect 430 454 433 456
rect 425 449 433 454
rect 435 454 443 458
rect 435 452 438 454
rect 440 452 443 454
rect 435 449 443 452
rect 379 446 381 448
rect 383 446 385 448
rect 379 444 385 446
rect 438 446 443 449
rect 445 446 450 458
rect 452 446 460 458
rect 510 457 515 458
rect 464 455 471 457
rect 464 453 466 455
rect 468 453 471 455
rect 464 451 471 453
rect 473 455 481 457
rect 473 453 476 455
rect 478 453 481 455
rect 473 451 481 453
rect 454 444 460 446
rect 454 442 456 444
rect 458 442 460 444
rect 454 440 460 442
rect 475 449 481 451
rect 483 449 488 457
rect 490 453 498 457
rect 490 451 493 453
rect 495 451 498 453
rect 490 449 498 451
rect 500 449 505 457
rect 507 453 515 457
rect 507 451 510 453
rect 512 451 515 453
rect 507 449 515 451
rect 517 456 524 458
rect 574 457 579 458
rect 517 454 520 456
rect 522 454 524 456
rect 517 452 524 454
rect 528 455 535 457
rect 528 453 530 455
rect 532 453 535 455
rect 517 449 522 452
rect 528 451 535 453
rect 537 455 545 457
rect 537 453 540 455
rect 542 453 545 455
rect 537 451 545 453
rect 539 449 545 451
rect 547 449 552 457
rect 554 453 562 457
rect 554 451 557 453
rect 559 451 562 453
rect 554 449 562 451
rect 564 449 569 457
rect 571 453 579 457
rect 571 451 574 453
rect 576 451 579 453
rect 571 449 579 451
rect 581 456 588 458
rect 638 457 643 458
rect 581 454 584 456
rect 586 454 588 456
rect 581 452 588 454
rect 592 455 599 457
rect 592 453 594 455
rect 596 453 599 455
rect 581 449 586 452
rect 592 451 599 453
rect 601 455 609 457
rect 601 453 604 455
rect 606 453 609 455
rect 601 451 609 453
rect 603 449 609 451
rect 611 449 616 457
rect 618 453 626 457
rect 618 451 621 453
rect 623 451 626 453
rect 618 449 626 451
rect 628 449 633 457
rect 635 453 643 457
rect 635 451 638 453
rect 640 451 643 453
rect 635 449 643 451
rect 645 456 652 458
rect 645 454 648 456
rect 650 454 652 456
rect 645 452 652 454
rect 645 449 650 452
rect 7 432 13 434
rect 7 430 9 432
rect 11 430 13 432
rect 7 428 13 430
rect 7 416 15 428
rect 17 416 22 428
rect 24 425 29 428
rect 89 432 96 434
rect 89 430 92 432
rect 94 430 96 432
rect 24 422 32 425
rect 24 420 27 422
rect 29 420 32 422
rect 24 416 32 420
rect 34 420 42 425
rect 34 418 37 420
rect 39 418 42 420
rect 34 416 42 418
rect 44 423 53 425
rect 89 424 96 430
rect 111 432 117 434
rect 111 430 113 432
rect 115 430 117 432
rect 111 428 117 430
rect 44 421 49 423
rect 51 421 53 423
rect 44 420 53 421
rect 71 422 78 424
rect 71 420 73 422
rect 75 420 78 422
rect 44 416 58 420
rect 53 411 58 416
rect 60 417 65 420
rect 71 418 78 420
rect 60 415 67 417
rect 60 413 63 415
rect 65 413 67 415
rect 73 413 78 418
rect 80 413 85 424
rect 87 422 96 424
rect 87 413 98 422
rect 100 420 107 422
rect 100 418 103 420
rect 105 418 107 420
rect 100 416 107 418
rect 111 416 119 428
rect 121 416 126 428
rect 128 425 133 428
rect 193 432 200 434
rect 193 430 196 432
rect 198 430 200 432
rect 128 422 136 425
rect 128 420 131 422
rect 133 420 136 422
rect 128 416 136 420
rect 138 420 146 425
rect 138 418 141 420
rect 143 418 146 420
rect 138 416 146 418
rect 148 423 157 425
rect 193 424 200 430
rect 215 428 221 430
rect 215 426 217 428
rect 219 426 221 428
rect 148 421 153 423
rect 155 421 157 423
rect 148 420 157 421
rect 175 422 182 424
rect 175 420 177 422
rect 179 420 182 422
rect 148 416 162 420
rect 100 413 105 416
rect 60 411 67 413
rect 157 411 162 416
rect 164 417 169 420
rect 175 418 182 420
rect 164 415 171 417
rect 164 413 167 415
rect 169 413 171 415
rect 177 413 182 418
rect 184 413 189 424
rect 191 422 200 424
rect 215 424 221 426
rect 234 428 240 430
rect 256 432 262 434
rect 256 430 258 432
rect 260 430 262 432
rect 256 428 262 430
rect 234 426 236 428
rect 238 426 240 428
rect 234 424 240 426
rect 191 413 202 422
rect 204 420 211 422
rect 204 418 207 420
rect 209 418 211 420
rect 204 416 211 418
rect 215 417 220 424
rect 236 420 240 424
rect 236 417 242 420
rect 204 413 209 416
rect 164 411 171 413
rect 215 411 222 417
rect 224 415 232 417
rect 224 413 227 415
rect 229 413 232 415
rect 224 411 232 413
rect 234 411 242 417
rect 244 417 249 420
rect 244 415 251 417
rect 256 416 264 428
rect 266 416 271 428
rect 273 425 278 428
rect 338 432 345 434
rect 338 430 341 432
rect 343 430 345 432
rect 273 422 281 425
rect 273 420 276 422
rect 278 420 281 422
rect 273 416 281 420
rect 283 420 291 425
rect 283 418 286 420
rect 288 418 291 420
rect 283 416 291 418
rect 293 423 302 425
rect 338 424 345 430
rect 360 428 366 430
rect 360 426 362 428
rect 364 426 366 428
rect 293 421 298 423
rect 300 421 302 423
rect 293 420 302 421
rect 320 422 327 424
rect 320 420 322 422
rect 324 420 327 422
rect 293 416 307 420
rect 244 413 247 415
rect 249 413 251 415
rect 244 411 251 413
rect 302 411 307 416
rect 309 417 314 420
rect 320 418 327 420
rect 309 415 316 417
rect 309 413 312 415
rect 314 413 316 415
rect 322 413 327 418
rect 329 413 334 424
rect 336 422 345 424
rect 360 424 366 426
rect 379 428 385 430
rect 379 426 381 428
rect 383 426 385 428
rect 379 424 385 426
rect 454 432 460 434
rect 454 430 456 432
rect 458 430 460 432
rect 454 428 460 430
rect 438 425 443 428
rect 336 413 347 422
rect 349 420 356 422
rect 349 418 352 420
rect 354 418 356 420
rect 349 416 356 418
rect 360 417 365 424
rect 381 420 385 424
rect 414 423 423 425
rect 414 421 416 423
rect 418 421 423 423
rect 414 420 423 421
rect 381 417 387 420
rect 349 413 354 416
rect 309 411 316 413
rect 360 411 367 417
rect 369 415 377 417
rect 369 413 372 415
rect 374 413 377 415
rect 369 411 377 413
rect 379 411 387 417
rect 389 417 394 420
rect 402 417 407 420
rect 389 415 396 417
rect 389 413 392 415
rect 394 413 396 415
rect 389 411 396 413
rect 400 415 407 417
rect 400 413 402 415
rect 404 413 407 415
rect 400 411 407 413
rect 409 416 423 420
rect 425 420 433 425
rect 425 418 428 420
rect 430 418 433 420
rect 425 416 433 418
rect 435 422 443 425
rect 435 420 438 422
rect 440 420 443 422
rect 435 416 443 420
rect 445 416 450 428
rect 452 416 460 428
rect 475 423 481 425
rect 464 421 471 423
rect 464 419 466 421
rect 468 419 471 421
rect 464 417 471 419
rect 473 421 481 423
rect 473 419 476 421
rect 478 419 481 421
rect 473 417 481 419
rect 483 417 488 425
rect 490 423 498 425
rect 490 421 493 423
rect 495 421 498 423
rect 490 417 498 421
rect 500 417 505 425
rect 507 423 515 425
rect 507 421 510 423
rect 512 421 515 423
rect 507 417 515 421
rect 409 411 414 416
rect 510 416 515 417
rect 517 422 522 425
rect 539 423 545 425
rect 517 420 524 422
rect 517 418 520 420
rect 522 418 524 420
rect 517 416 524 418
rect 528 421 535 423
rect 528 419 530 421
rect 532 419 535 421
rect 528 417 535 419
rect 537 421 545 423
rect 537 419 540 421
rect 542 419 545 421
rect 537 417 545 419
rect 547 417 552 425
rect 554 423 562 425
rect 554 421 557 423
rect 559 421 562 423
rect 554 417 562 421
rect 564 417 569 425
rect 571 423 579 425
rect 571 421 574 423
rect 576 421 579 423
rect 571 417 579 421
rect 574 416 579 417
rect 581 422 586 425
rect 603 423 609 425
rect 581 420 588 422
rect 581 418 584 420
rect 586 418 588 420
rect 581 416 588 418
rect 592 421 599 423
rect 592 419 594 421
rect 596 419 599 421
rect 592 417 599 419
rect 601 421 609 423
rect 601 419 604 421
rect 606 419 609 421
rect 601 417 609 419
rect 611 417 616 425
rect 618 423 626 425
rect 618 421 621 423
rect 623 421 626 423
rect 618 417 626 421
rect 628 417 633 425
rect 635 423 643 425
rect 635 421 638 423
rect 640 421 643 423
rect 635 417 643 421
rect 638 416 643 417
rect 645 422 650 425
rect 645 420 652 422
rect 645 418 648 420
rect 650 418 652 420
rect 645 416 652 418
rect 7 317 14 319
rect 7 315 9 317
rect 11 315 14 317
rect 7 313 14 315
rect 9 310 14 313
rect 16 313 24 319
rect 26 317 34 319
rect 26 315 29 317
rect 31 315 34 317
rect 26 313 34 315
rect 36 313 43 319
rect 87 317 94 319
rect 49 314 54 317
rect 16 310 22 313
rect 18 306 22 310
rect 38 306 43 313
rect 47 312 54 314
rect 47 310 49 312
rect 51 310 54 312
rect 47 308 54 310
rect 56 308 67 317
rect 18 304 24 306
rect 18 302 20 304
rect 22 302 24 304
rect 18 300 24 302
rect 37 304 43 306
rect 58 306 67 308
rect 69 306 74 317
rect 76 312 81 317
rect 87 315 89 317
rect 91 315 94 317
rect 87 313 94 315
rect 76 310 83 312
rect 89 310 94 313
rect 96 314 101 319
rect 191 317 198 319
rect 153 314 158 317
rect 96 310 110 314
rect 76 308 79 310
rect 81 308 83 310
rect 76 306 83 308
rect 101 309 110 310
rect 101 307 103 309
rect 105 307 110 309
rect 37 302 39 304
rect 41 302 43 304
rect 37 300 43 302
rect 58 300 65 306
rect 101 305 110 307
rect 112 312 120 314
rect 112 310 115 312
rect 117 310 120 312
rect 112 305 120 310
rect 122 310 130 314
rect 122 308 125 310
rect 127 308 130 310
rect 122 305 130 308
rect 58 298 60 300
rect 62 298 65 300
rect 58 296 65 298
rect 125 302 130 305
rect 132 302 137 314
rect 139 302 147 314
rect 151 312 158 314
rect 151 310 153 312
rect 155 310 158 312
rect 151 308 158 310
rect 160 308 171 317
rect 162 306 171 308
rect 173 306 178 317
rect 180 312 185 317
rect 191 315 193 317
rect 195 315 198 317
rect 191 313 198 315
rect 180 310 187 312
rect 193 310 198 313
rect 200 314 205 319
rect 302 314 307 319
rect 200 310 214 314
rect 180 308 183 310
rect 185 308 187 310
rect 180 306 187 308
rect 205 309 214 310
rect 205 307 207 309
rect 209 307 214 309
rect 141 300 147 302
rect 141 298 143 300
rect 145 298 147 300
rect 141 296 147 298
rect 162 300 169 306
rect 205 305 214 307
rect 216 312 224 314
rect 216 310 219 312
rect 221 310 224 312
rect 216 305 224 310
rect 226 310 234 314
rect 226 308 229 310
rect 231 308 234 310
rect 226 305 234 308
rect 162 298 164 300
rect 166 298 169 300
rect 162 296 169 298
rect 229 302 234 305
rect 236 302 241 314
rect 243 302 251 314
rect 245 300 251 302
rect 245 298 247 300
rect 249 298 251 300
rect 245 296 251 298
rect 256 302 264 314
rect 266 302 271 314
rect 273 310 281 314
rect 273 308 276 310
rect 278 308 281 310
rect 273 305 281 308
rect 283 312 291 314
rect 283 310 286 312
rect 288 310 291 312
rect 283 305 291 310
rect 293 310 307 314
rect 309 317 316 319
rect 309 315 312 317
rect 314 315 316 317
rect 309 313 316 315
rect 309 310 314 313
rect 322 312 327 317
rect 320 310 327 312
rect 293 309 302 310
rect 293 307 298 309
rect 300 307 302 309
rect 293 305 302 307
rect 320 308 322 310
rect 324 308 327 310
rect 320 306 327 308
rect 329 306 334 317
rect 336 308 347 317
rect 349 314 354 317
rect 349 312 356 314
rect 349 310 352 312
rect 354 310 356 312
rect 349 308 356 310
rect 360 313 367 319
rect 369 317 377 319
rect 369 315 372 317
rect 374 315 377 317
rect 369 313 377 315
rect 379 313 387 319
rect 336 306 345 308
rect 273 302 278 305
rect 256 300 262 302
rect 256 298 258 300
rect 260 298 262 300
rect 256 296 262 298
rect 338 300 345 306
rect 360 306 365 313
rect 381 310 387 313
rect 389 317 396 319
rect 389 315 392 317
rect 394 315 396 317
rect 389 313 396 315
rect 400 317 407 319
rect 400 315 402 317
rect 404 315 407 317
rect 400 313 407 315
rect 389 310 394 313
rect 402 310 407 313
rect 409 314 414 319
rect 409 310 423 314
rect 381 306 385 310
rect 360 304 366 306
rect 360 302 362 304
rect 364 302 366 304
rect 338 298 341 300
rect 343 298 345 300
rect 338 296 345 298
rect 360 300 366 302
rect 379 304 385 306
rect 414 309 423 310
rect 414 307 416 309
rect 418 307 423 309
rect 414 305 423 307
rect 425 312 433 314
rect 425 310 428 312
rect 430 310 433 312
rect 425 305 433 310
rect 435 310 443 314
rect 435 308 438 310
rect 440 308 443 310
rect 435 305 443 308
rect 379 302 381 304
rect 383 302 385 304
rect 379 300 385 302
rect 438 302 443 305
rect 445 302 450 314
rect 452 302 460 314
rect 510 313 515 314
rect 464 311 471 313
rect 464 309 466 311
rect 468 309 471 311
rect 464 307 471 309
rect 473 311 481 313
rect 473 309 476 311
rect 478 309 481 311
rect 473 307 481 309
rect 454 300 460 302
rect 454 298 456 300
rect 458 298 460 300
rect 454 296 460 298
rect 475 305 481 307
rect 483 305 488 313
rect 490 309 498 313
rect 490 307 493 309
rect 495 307 498 309
rect 490 305 498 307
rect 500 305 505 313
rect 507 309 515 313
rect 507 307 510 309
rect 512 307 515 309
rect 507 305 515 307
rect 517 312 524 314
rect 574 313 579 314
rect 517 310 520 312
rect 522 310 524 312
rect 517 308 524 310
rect 528 311 535 313
rect 528 309 530 311
rect 532 309 535 311
rect 517 305 522 308
rect 528 307 535 309
rect 537 311 545 313
rect 537 309 540 311
rect 542 309 545 311
rect 537 307 545 309
rect 539 305 545 307
rect 547 305 552 313
rect 554 309 562 313
rect 554 307 557 309
rect 559 307 562 309
rect 554 305 562 307
rect 564 305 569 313
rect 571 309 579 313
rect 571 307 574 309
rect 576 307 579 309
rect 571 305 579 307
rect 581 312 588 314
rect 638 313 643 314
rect 581 310 584 312
rect 586 310 588 312
rect 581 308 588 310
rect 592 311 599 313
rect 592 309 594 311
rect 596 309 599 311
rect 581 305 586 308
rect 592 307 599 309
rect 601 311 609 313
rect 601 309 604 311
rect 606 309 609 311
rect 601 307 609 309
rect 603 305 609 307
rect 611 305 616 313
rect 618 309 626 313
rect 618 307 621 309
rect 623 307 626 309
rect 618 305 626 307
rect 628 305 633 313
rect 635 309 643 313
rect 635 307 638 309
rect 640 307 643 309
rect 635 305 643 307
rect 645 312 652 314
rect 645 310 648 312
rect 650 310 652 312
rect 645 308 652 310
rect 645 305 650 308
rect 7 288 13 290
rect 7 286 9 288
rect 11 286 13 288
rect 7 284 13 286
rect 7 272 15 284
rect 17 272 22 284
rect 24 281 29 284
rect 89 288 96 290
rect 89 286 92 288
rect 94 286 96 288
rect 24 278 32 281
rect 24 276 27 278
rect 29 276 32 278
rect 24 272 32 276
rect 34 276 42 281
rect 34 274 37 276
rect 39 274 42 276
rect 34 272 42 274
rect 44 279 53 281
rect 89 280 96 286
rect 111 288 117 290
rect 111 286 113 288
rect 115 286 117 288
rect 111 284 117 286
rect 44 277 49 279
rect 51 277 53 279
rect 44 276 53 277
rect 71 278 78 280
rect 71 276 73 278
rect 75 276 78 278
rect 44 272 58 276
rect 53 267 58 272
rect 60 273 65 276
rect 71 274 78 276
rect 60 271 67 273
rect 60 269 63 271
rect 65 269 67 271
rect 73 269 78 274
rect 80 269 85 280
rect 87 278 96 280
rect 87 269 98 278
rect 100 276 107 278
rect 100 274 103 276
rect 105 274 107 276
rect 100 272 107 274
rect 111 272 119 284
rect 121 272 126 284
rect 128 281 133 284
rect 193 288 200 290
rect 193 286 196 288
rect 198 286 200 288
rect 128 278 136 281
rect 128 276 131 278
rect 133 276 136 278
rect 128 272 136 276
rect 138 276 146 281
rect 138 274 141 276
rect 143 274 146 276
rect 138 272 146 274
rect 148 279 157 281
rect 193 280 200 286
rect 215 284 221 286
rect 215 282 217 284
rect 219 282 221 284
rect 148 277 153 279
rect 155 277 157 279
rect 148 276 157 277
rect 175 278 182 280
rect 175 276 177 278
rect 179 276 182 278
rect 148 272 162 276
rect 100 269 105 272
rect 60 267 67 269
rect 157 267 162 272
rect 164 273 169 276
rect 175 274 182 276
rect 164 271 171 273
rect 164 269 167 271
rect 169 269 171 271
rect 177 269 182 274
rect 184 269 189 280
rect 191 278 200 280
rect 215 280 221 282
rect 234 284 240 286
rect 256 288 262 290
rect 256 286 258 288
rect 260 286 262 288
rect 256 284 262 286
rect 234 282 236 284
rect 238 282 240 284
rect 234 280 240 282
rect 191 269 202 278
rect 204 276 211 278
rect 204 274 207 276
rect 209 274 211 276
rect 204 272 211 274
rect 215 273 220 280
rect 236 276 240 280
rect 236 273 242 276
rect 204 269 209 272
rect 164 267 171 269
rect 215 267 222 273
rect 224 271 232 273
rect 224 269 227 271
rect 229 269 232 271
rect 224 267 232 269
rect 234 267 242 273
rect 244 273 249 276
rect 244 271 251 273
rect 256 272 264 284
rect 266 272 271 284
rect 273 281 278 284
rect 338 288 345 290
rect 338 286 341 288
rect 343 286 345 288
rect 273 278 281 281
rect 273 276 276 278
rect 278 276 281 278
rect 273 272 281 276
rect 283 276 291 281
rect 283 274 286 276
rect 288 274 291 276
rect 283 272 291 274
rect 293 279 302 281
rect 338 280 345 286
rect 360 284 366 286
rect 360 282 362 284
rect 364 282 366 284
rect 293 277 298 279
rect 300 277 302 279
rect 293 276 302 277
rect 320 278 327 280
rect 320 276 322 278
rect 324 276 327 278
rect 293 272 307 276
rect 244 269 247 271
rect 249 269 251 271
rect 244 267 251 269
rect 302 267 307 272
rect 309 273 314 276
rect 320 274 327 276
rect 309 271 316 273
rect 309 269 312 271
rect 314 269 316 271
rect 322 269 327 274
rect 329 269 334 280
rect 336 278 345 280
rect 360 280 366 282
rect 379 284 385 286
rect 379 282 381 284
rect 383 282 385 284
rect 379 280 385 282
rect 454 288 460 290
rect 454 286 456 288
rect 458 286 460 288
rect 454 284 460 286
rect 438 281 443 284
rect 336 269 347 278
rect 349 276 356 278
rect 349 274 352 276
rect 354 274 356 276
rect 349 272 356 274
rect 360 273 365 280
rect 381 276 385 280
rect 414 279 423 281
rect 414 277 416 279
rect 418 277 423 279
rect 414 276 423 277
rect 381 273 387 276
rect 349 269 354 272
rect 309 267 316 269
rect 360 267 367 273
rect 369 271 377 273
rect 369 269 372 271
rect 374 269 377 271
rect 369 267 377 269
rect 379 267 387 273
rect 389 273 394 276
rect 402 273 407 276
rect 389 271 396 273
rect 389 269 392 271
rect 394 269 396 271
rect 389 267 396 269
rect 400 271 407 273
rect 400 269 402 271
rect 404 269 407 271
rect 400 267 407 269
rect 409 272 423 276
rect 425 276 433 281
rect 425 274 428 276
rect 430 274 433 276
rect 425 272 433 274
rect 435 278 443 281
rect 435 276 438 278
rect 440 276 443 278
rect 435 272 443 276
rect 445 272 450 284
rect 452 272 460 284
rect 475 279 481 281
rect 464 277 471 279
rect 464 275 466 277
rect 468 275 471 277
rect 464 273 471 275
rect 473 277 481 279
rect 473 275 476 277
rect 478 275 481 277
rect 473 273 481 275
rect 483 273 488 281
rect 490 279 498 281
rect 490 277 493 279
rect 495 277 498 279
rect 490 273 498 277
rect 500 273 505 281
rect 507 279 515 281
rect 507 277 510 279
rect 512 277 515 279
rect 507 273 515 277
rect 409 267 414 272
rect 510 272 515 273
rect 517 278 522 281
rect 539 279 545 281
rect 517 276 524 278
rect 517 274 520 276
rect 522 274 524 276
rect 517 272 524 274
rect 528 277 535 279
rect 528 275 530 277
rect 532 275 535 277
rect 528 273 535 275
rect 537 277 545 279
rect 537 275 540 277
rect 542 275 545 277
rect 537 273 545 275
rect 547 273 552 281
rect 554 279 562 281
rect 554 277 557 279
rect 559 277 562 279
rect 554 273 562 277
rect 564 273 569 281
rect 571 279 579 281
rect 571 277 574 279
rect 576 277 579 279
rect 571 273 579 277
rect 574 272 579 273
rect 581 278 586 281
rect 603 279 609 281
rect 581 276 588 278
rect 581 274 584 276
rect 586 274 588 276
rect 581 272 588 274
rect 592 277 599 279
rect 592 275 594 277
rect 596 275 599 277
rect 592 273 599 275
rect 601 277 609 279
rect 601 275 604 277
rect 606 275 609 277
rect 601 273 609 275
rect 611 273 616 281
rect 618 279 626 281
rect 618 277 621 279
rect 623 277 626 279
rect 618 273 626 277
rect 628 273 633 281
rect 635 279 643 281
rect 635 277 638 279
rect 640 277 643 279
rect 635 273 643 277
rect 638 272 643 273
rect 645 278 650 281
rect 645 276 652 278
rect 645 274 648 276
rect 650 274 652 276
rect 645 272 652 274
rect 7 173 14 175
rect 7 171 9 173
rect 11 171 14 173
rect 7 169 14 171
rect 9 166 14 169
rect 16 169 24 175
rect 26 173 34 175
rect 26 171 29 173
rect 31 171 34 173
rect 26 169 34 171
rect 36 169 43 175
rect 87 173 94 175
rect 49 170 54 173
rect 16 166 22 169
rect 18 162 22 166
rect 38 162 43 169
rect 47 168 54 170
rect 47 166 49 168
rect 51 166 54 168
rect 47 164 54 166
rect 56 164 67 173
rect 18 160 24 162
rect 18 158 20 160
rect 22 158 24 160
rect 18 156 24 158
rect 37 160 43 162
rect 58 162 67 164
rect 69 162 74 173
rect 76 168 81 173
rect 87 171 89 173
rect 91 171 94 173
rect 87 169 94 171
rect 76 166 83 168
rect 89 166 94 169
rect 96 170 101 175
rect 191 173 198 175
rect 153 170 158 173
rect 96 166 110 170
rect 76 164 79 166
rect 81 164 83 166
rect 76 162 83 164
rect 101 165 110 166
rect 101 163 103 165
rect 105 163 110 165
rect 37 158 39 160
rect 41 158 43 160
rect 37 156 43 158
rect 58 156 65 162
rect 101 161 110 163
rect 112 168 120 170
rect 112 166 115 168
rect 117 166 120 168
rect 112 161 120 166
rect 122 166 130 170
rect 122 164 125 166
rect 127 164 130 166
rect 122 161 130 164
rect 58 154 60 156
rect 62 154 65 156
rect 58 152 65 154
rect 125 158 130 161
rect 132 158 137 170
rect 139 158 147 170
rect 151 168 158 170
rect 151 166 153 168
rect 155 166 158 168
rect 151 164 158 166
rect 160 164 171 173
rect 162 162 171 164
rect 173 162 178 173
rect 180 168 185 173
rect 191 171 193 173
rect 195 171 198 173
rect 191 169 198 171
rect 180 166 187 168
rect 193 166 198 169
rect 200 170 205 175
rect 302 170 307 175
rect 200 166 214 170
rect 180 164 183 166
rect 185 164 187 166
rect 180 162 187 164
rect 205 165 214 166
rect 205 163 207 165
rect 209 163 214 165
rect 141 156 147 158
rect 141 154 143 156
rect 145 154 147 156
rect 141 152 147 154
rect 162 156 169 162
rect 205 161 214 163
rect 216 168 224 170
rect 216 166 219 168
rect 221 166 224 168
rect 216 161 224 166
rect 226 166 234 170
rect 226 164 229 166
rect 231 164 234 166
rect 226 161 234 164
rect 162 154 164 156
rect 166 154 169 156
rect 162 152 169 154
rect 229 158 234 161
rect 236 158 241 170
rect 243 158 251 170
rect 245 156 251 158
rect 245 154 247 156
rect 249 154 251 156
rect 245 152 251 154
rect 256 158 264 170
rect 266 158 271 170
rect 273 166 281 170
rect 273 164 276 166
rect 278 164 281 166
rect 273 161 281 164
rect 283 168 291 170
rect 283 166 286 168
rect 288 166 291 168
rect 283 161 291 166
rect 293 166 307 170
rect 309 173 316 175
rect 309 171 312 173
rect 314 171 316 173
rect 309 169 316 171
rect 309 166 314 169
rect 322 168 327 173
rect 320 166 327 168
rect 293 165 302 166
rect 293 163 298 165
rect 300 163 302 165
rect 293 161 302 163
rect 320 164 322 166
rect 324 164 327 166
rect 320 162 327 164
rect 329 162 334 173
rect 336 164 347 173
rect 349 170 354 173
rect 349 168 356 170
rect 349 166 352 168
rect 354 166 356 168
rect 349 164 356 166
rect 360 169 367 175
rect 369 173 377 175
rect 369 171 372 173
rect 374 171 377 173
rect 369 169 377 171
rect 379 169 387 175
rect 336 162 345 164
rect 273 158 278 161
rect 256 156 262 158
rect 256 154 258 156
rect 260 154 262 156
rect 256 152 262 154
rect 338 156 345 162
rect 360 162 365 169
rect 381 166 387 169
rect 389 173 396 175
rect 389 171 392 173
rect 394 171 396 173
rect 389 169 396 171
rect 400 173 407 175
rect 400 171 402 173
rect 404 171 407 173
rect 400 169 407 171
rect 389 166 394 169
rect 402 166 407 169
rect 409 170 414 175
rect 409 166 423 170
rect 381 162 385 166
rect 360 160 366 162
rect 360 158 362 160
rect 364 158 366 160
rect 338 154 341 156
rect 343 154 345 156
rect 338 152 345 154
rect 360 156 366 158
rect 379 160 385 162
rect 414 165 423 166
rect 414 163 416 165
rect 418 163 423 165
rect 414 161 423 163
rect 425 168 433 170
rect 425 166 428 168
rect 430 166 433 168
rect 425 161 433 166
rect 435 166 443 170
rect 435 164 438 166
rect 440 164 443 166
rect 435 161 443 164
rect 379 158 381 160
rect 383 158 385 160
rect 379 156 385 158
rect 438 158 443 161
rect 445 158 450 170
rect 452 158 460 170
rect 510 169 515 170
rect 464 167 471 169
rect 464 165 466 167
rect 468 165 471 167
rect 464 163 471 165
rect 473 167 481 169
rect 473 165 476 167
rect 478 165 481 167
rect 473 163 481 165
rect 454 156 460 158
rect 454 154 456 156
rect 458 154 460 156
rect 454 152 460 154
rect 475 161 481 163
rect 483 161 488 169
rect 490 165 498 169
rect 490 163 493 165
rect 495 163 498 165
rect 490 161 498 163
rect 500 161 505 169
rect 507 165 515 169
rect 507 163 510 165
rect 512 163 515 165
rect 507 161 515 163
rect 517 168 524 170
rect 574 169 579 170
rect 517 166 520 168
rect 522 166 524 168
rect 517 164 524 166
rect 528 167 535 169
rect 528 165 530 167
rect 532 165 535 167
rect 517 161 522 164
rect 528 163 535 165
rect 537 167 545 169
rect 537 165 540 167
rect 542 165 545 167
rect 537 163 545 165
rect 539 161 545 163
rect 547 161 552 169
rect 554 165 562 169
rect 554 163 557 165
rect 559 163 562 165
rect 554 161 562 163
rect 564 161 569 169
rect 571 165 579 169
rect 571 163 574 165
rect 576 163 579 165
rect 571 161 579 163
rect 581 168 588 170
rect 638 169 643 170
rect 581 166 584 168
rect 586 166 588 168
rect 581 164 588 166
rect 592 167 599 169
rect 592 165 594 167
rect 596 165 599 167
rect 581 161 586 164
rect 592 163 599 165
rect 601 167 609 169
rect 601 165 604 167
rect 606 165 609 167
rect 601 163 609 165
rect 603 161 609 163
rect 611 161 616 169
rect 618 165 626 169
rect 618 163 621 165
rect 623 163 626 165
rect 618 161 626 163
rect 628 161 633 169
rect 635 165 643 169
rect 635 163 638 165
rect 640 163 643 165
rect 635 161 643 163
rect 645 168 652 170
rect 645 166 648 168
rect 650 166 652 168
rect 645 164 652 166
rect 645 161 650 164
rect 7 144 13 146
rect 7 142 9 144
rect 11 142 13 144
rect 7 140 13 142
rect 7 128 15 140
rect 17 128 22 140
rect 24 137 29 140
rect 89 144 96 146
rect 89 142 92 144
rect 94 142 96 144
rect 24 134 32 137
rect 24 132 27 134
rect 29 132 32 134
rect 24 128 32 132
rect 34 132 42 137
rect 34 130 37 132
rect 39 130 42 132
rect 34 128 42 130
rect 44 135 53 137
rect 89 136 96 142
rect 111 144 117 146
rect 111 142 113 144
rect 115 142 117 144
rect 111 140 117 142
rect 44 133 49 135
rect 51 133 53 135
rect 44 132 53 133
rect 71 134 78 136
rect 71 132 73 134
rect 75 132 78 134
rect 44 128 58 132
rect 53 123 58 128
rect 60 129 65 132
rect 71 130 78 132
rect 60 127 67 129
rect 60 125 63 127
rect 65 125 67 127
rect 73 125 78 130
rect 80 125 85 136
rect 87 134 96 136
rect 87 125 98 134
rect 100 132 107 134
rect 100 130 103 132
rect 105 130 107 132
rect 100 128 107 130
rect 111 128 119 140
rect 121 128 126 140
rect 128 137 133 140
rect 193 144 200 146
rect 193 142 196 144
rect 198 142 200 144
rect 128 134 136 137
rect 128 132 131 134
rect 133 132 136 134
rect 128 128 136 132
rect 138 132 146 137
rect 138 130 141 132
rect 143 130 146 132
rect 138 128 146 130
rect 148 135 157 137
rect 193 136 200 142
rect 215 140 221 142
rect 215 138 217 140
rect 219 138 221 140
rect 148 133 153 135
rect 155 133 157 135
rect 148 132 157 133
rect 175 134 182 136
rect 175 132 177 134
rect 179 132 182 134
rect 148 128 162 132
rect 100 125 105 128
rect 60 123 67 125
rect 157 123 162 128
rect 164 129 169 132
rect 175 130 182 132
rect 164 127 171 129
rect 164 125 167 127
rect 169 125 171 127
rect 177 125 182 130
rect 184 125 189 136
rect 191 134 200 136
rect 215 136 221 138
rect 234 140 240 142
rect 256 144 262 146
rect 256 142 258 144
rect 260 142 262 144
rect 256 140 262 142
rect 234 138 236 140
rect 238 138 240 140
rect 234 136 240 138
rect 191 125 202 134
rect 204 132 211 134
rect 204 130 207 132
rect 209 130 211 132
rect 204 128 211 130
rect 215 129 220 136
rect 236 132 240 136
rect 236 129 242 132
rect 204 125 209 128
rect 164 123 171 125
rect 215 123 222 129
rect 224 127 232 129
rect 224 125 227 127
rect 229 125 232 127
rect 224 123 232 125
rect 234 123 242 129
rect 244 129 249 132
rect 244 127 251 129
rect 256 128 264 140
rect 266 128 271 140
rect 273 137 278 140
rect 338 144 345 146
rect 338 142 341 144
rect 343 142 345 144
rect 273 134 281 137
rect 273 132 276 134
rect 278 132 281 134
rect 273 128 281 132
rect 283 132 291 137
rect 283 130 286 132
rect 288 130 291 132
rect 283 128 291 130
rect 293 135 302 137
rect 338 136 345 142
rect 360 140 366 142
rect 360 138 362 140
rect 364 138 366 140
rect 293 133 298 135
rect 300 133 302 135
rect 293 132 302 133
rect 320 134 327 136
rect 320 132 322 134
rect 324 132 327 134
rect 293 128 307 132
rect 244 125 247 127
rect 249 125 251 127
rect 244 123 251 125
rect 302 123 307 128
rect 309 129 314 132
rect 320 130 327 132
rect 309 127 316 129
rect 309 125 312 127
rect 314 125 316 127
rect 322 125 327 130
rect 329 125 334 136
rect 336 134 345 136
rect 360 136 366 138
rect 379 140 385 142
rect 379 138 381 140
rect 383 138 385 140
rect 379 136 385 138
rect 454 144 460 146
rect 454 142 456 144
rect 458 142 460 144
rect 454 140 460 142
rect 438 137 443 140
rect 336 125 347 134
rect 349 132 356 134
rect 349 130 352 132
rect 354 130 356 132
rect 349 128 356 130
rect 360 129 365 136
rect 381 132 385 136
rect 414 135 423 137
rect 414 133 416 135
rect 418 133 423 135
rect 414 132 423 133
rect 381 129 387 132
rect 349 125 354 128
rect 309 123 316 125
rect 360 123 367 129
rect 369 127 377 129
rect 369 125 372 127
rect 374 125 377 127
rect 369 123 377 125
rect 379 123 387 129
rect 389 129 394 132
rect 402 129 407 132
rect 389 127 396 129
rect 389 125 392 127
rect 394 125 396 127
rect 389 123 396 125
rect 400 127 407 129
rect 400 125 402 127
rect 404 125 407 127
rect 400 123 407 125
rect 409 128 423 132
rect 425 132 433 137
rect 425 130 428 132
rect 430 130 433 132
rect 425 128 433 130
rect 435 134 443 137
rect 435 132 438 134
rect 440 132 443 134
rect 435 128 443 132
rect 445 128 450 140
rect 452 128 460 140
rect 475 135 481 137
rect 464 133 471 135
rect 464 131 466 133
rect 468 131 471 133
rect 464 129 471 131
rect 473 133 481 135
rect 473 131 476 133
rect 478 131 481 133
rect 473 129 481 131
rect 483 129 488 137
rect 490 135 498 137
rect 490 133 493 135
rect 495 133 498 135
rect 490 129 498 133
rect 500 129 505 137
rect 507 135 515 137
rect 507 133 510 135
rect 512 133 515 135
rect 507 129 515 133
rect 409 123 414 128
rect 510 128 515 129
rect 517 134 522 137
rect 539 135 545 137
rect 517 132 524 134
rect 517 130 520 132
rect 522 130 524 132
rect 517 128 524 130
rect 528 133 535 135
rect 528 131 530 133
rect 532 131 535 133
rect 528 129 535 131
rect 537 133 545 135
rect 537 131 540 133
rect 542 131 545 133
rect 537 129 545 131
rect 547 129 552 137
rect 554 135 562 137
rect 554 133 557 135
rect 559 133 562 135
rect 554 129 562 133
rect 564 129 569 137
rect 571 135 579 137
rect 571 133 574 135
rect 576 133 579 135
rect 571 129 579 133
rect 574 128 579 129
rect 581 134 586 137
rect 603 135 609 137
rect 581 132 588 134
rect 581 130 584 132
rect 586 130 588 132
rect 581 128 588 130
rect 592 133 599 135
rect 592 131 594 133
rect 596 131 599 133
rect 592 129 599 131
rect 601 133 609 135
rect 601 131 604 133
rect 606 131 609 133
rect 601 129 609 131
rect 611 129 616 137
rect 618 135 626 137
rect 618 133 621 135
rect 623 133 626 135
rect 618 129 626 133
rect 628 129 633 137
rect 635 135 643 137
rect 635 133 638 135
rect 640 133 643 135
rect 635 129 643 133
rect 638 128 643 129
rect 645 134 650 137
rect 645 132 652 134
rect 645 130 648 132
rect 650 130 652 132
rect 645 128 652 130
rect 7 29 14 31
rect 7 27 9 29
rect 11 27 14 29
rect 7 25 14 27
rect 9 22 14 25
rect 16 25 24 31
rect 26 29 34 31
rect 26 27 29 29
rect 31 27 34 29
rect 26 25 34 27
rect 36 25 43 31
rect 87 29 94 31
rect 49 26 54 29
rect 16 22 22 25
rect 18 18 22 22
rect 38 18 43 25
rect 47 24 54 26
rect 47 22 49 24
rect 51 22 54 24
rect 47 20 54 22
rect 56 20 67 29
rect 18 16 24 18
rect 18 14 20 16
rect 22 14 24 16
rect 18 12 24 14
rect 37 16 43 18
rect 58 18 67 20
rect 69 18 74 29
rect 76 24 81 29
rect 87 27 89 29
rect 91 27 94 29
rect 87 25 94 27
rect 76 22 83 24
rect 89 22 94 25
rect 96 26 101 31
rect 191 29 198 31
rect 153 26 158 29
rect 96 22 110 26
rect 76 20 79 22
rect 81 20 83 22
rect 76 18 83 20
rect 101 21 110 22
rect 101 19 103 21
rect 105 19 110 21
rect 37 14 39 16
rect 41 14 43 16
rect 37 12 43 14
rect 58 12 65 18
rect 101 17 110 19
rect 112 24 120 26
rect 112 22 115 24
rect 117 22 120 24
rect 112 17 120 22
rect 122 22 130 26
rect 122 20 125 22
rect 127 20 130 22
rect 122 17 130 20
rect 58 10 60 12
rect 62 10 65 12
rect 58 8 65 10
rect 125 14 130 17
rect 132 14 137 26
rect 139 14 147 26
rect 151 24 158 26
rect 151 22 153 24
rect 155 22 158 24
rect 151 20 158 22
rect 160 20 171 29
rect 162 18 171 20
rect 173 18 178 29
rect 180 24 185 29
rect 191 27 193 29
rect 195 27 198 29
rect 191 25 198 27
rect 180 22 187 24
rect 193 22 198 25
rect 200 26 205 31
rect 302 26 307 31
rect 200 22 214 26
rect 180 20 183 22
rect 185 20 187 22
rect 180 18 187 20
rect 205 21 214 22
rect 205 19 207 21
rect 209 19 214 21
rect 141 12 147 14
rect 141 10 143 12
rect 145 10 147 12
rect 141 8 147 10
rect 162 12 169 18
rect 205 17 214 19
rect 216 24 224 26
rect 216 22 219 24
rect 221 22 224 24
rect 216 17 224 22
rect 226 22 234 26
rect 226 20 229 22
rect 231 20 234 22
rect 226 17 234 20
rect 162 10 164 12
rect 166 10 169 12
rect 162 8 169 10
rect 229 14 234 17
rect 236 14 241 26
rect 243 14 251 26
rect 245 12 251 14
rect 245 10 247 12
rect 249 10 251 12
rect 245 8 251 10
rect 256 14 264 26
rect 266 14 271 26
rect 273 22 281 26
rect 273 20 276 22
rect 278 20 281 22
rect 273 17 281 20
rect 283 24 291 26
rect 283 22 286 24
rect 288 22 291 24
rect 283 17 291 22
rect 293 22 307 26
rect 309 29 316 31
rect 309 27 312 29
rect 314 27 316 29
rect 309 25 316 27
rect 309 22 314 25
rect 322 24 327 29
rect 320 22 327 24
rect 293 21 302 22
rect 293 19 298 21
rect 300 19 302 21
rect 293 17 302 19
rect 320 20 322 22
rect 324 20 327 22
rect 320 18 327 20
rect 329 18 334 29
rect 336 20 347 29
rect 349 26 354 29
rect 349 24 356 26
rect 349 22 352 24
rect 354 22 356 24
rect 349 20 356 22
rect 360 25 367 31
rect 369 29 377 31
rect 369 27 372 29
rect 374 27 377 29
rect 369 25 377 27
rect 379 25 387 31
rect 336 18 345 20
rect 273 14 278 17
rect 256 12 262 14
rect 256 10 258 12
rect 260 10 262 12
rect 256 8 262 10
rect 338 12 345 18
rect 360 18 365 25
rect 381 22 387 25
rect 389 29 396 31
rect 389 27 392 29
rect 394 27 396 29
rect 389 25 396 27
rect 400 29 407 31
rect 400 27 402 29
rect 404 27 407 29
rect 400 25 407 27
rect 389 22 394 25
rect 402 22 407 25
rect 409 26 414 31
rect 409 22 423 26
rect 381 18 385 22
rect 360 16 366 18
rect 360 14 362 16
rect 364 14 366 16
rect 338 10 341 12
rect 343 10 345 12
rect 338 8 345 10
rect 360 12 366 14
rect 379 16 385 18
rect 414 21 423 22
rect 414 19 416 21
rect 418 19 423 21
rect 414 17 423 19
rect 425 24 433 26
rect 425 22 428 24
rect 430 22 433 24
rect 425 17 433 22
rect 435 22 443 26
rect 435 20 438 22
rect 440 20 443 22
rect 435 17 443 20
rect 379 14 381 16
rect 383 14 385 16
rect 379 12 385 14
rect 438 14 443 17
rect 445 14 450 26
rect 452 14 460 26
rect 510 25 515 26
rect 464 23 471 25
rect 464 21 466 23
rect 468 21 471 23
rect 464 19 471 21
rect 473 23 481 25
rect 473 21 476 23
rect 478 21 481 23
rect 473 19 481 21
rect 454 12 460 14
rect 454 10 456 12
rect 458 10 460 12
rect 454 8 460 10
rect 475 17 481 19
rect 483 17 488 25
rect 490 21 498 25
rect 490 19 493 21
rect 495 19 498 21
rect 490 17 498 19
rect 500 17 505 25
rect 507 21 515 25
rect 507 19 510 21
rect 512 19 515 21
rect 507 17 515 19
rect 517 24 524 26
rect 574 25 579 26
rect 517 22 520 24
rect 522 22 524 24
rect 517 20 524 22
rect 528 23 535 25
rect 528 21 530 23
rect 532 21 535 23
rect 517 17 522 20
rect 528 19 535 21
rect 537 23 545 25
rect 537 21 540 23
rect 542 21 545 23
rect 537 19 545 21
rect 539 17 545 19
rect 547 17 552 25
rect 554 21 562 25
rect 554 19 557 21
rect 559 19 562 21
rect 554 17 562 19
rect 564 17 569 25
rect 571 21 579 25
rect 571 19 574 21
rect 576 19 579 21
rect 571 17 579 19
rect 581 24 588 26
rect 638 25 643 26
rect 581 22 584 24
rect 586 22 588 24
rect 581 20 588 22
rect 592 23 599 25
rect 592 21 594 23
rect 596 21 599 23
rect 581 17 586 20
rect 592 19 599 21
rect 601 23 609 25
rect 601 21 604 23
rect 606 21 609 23
rect 601 19 609 21
rect 603 17 609 19
rect 611 17 616 25
rect 618 21 626 25
rect 618 19 621 21
rect 623 19 626 21
rect 618 17 626 19
rect 628 17 633 25
rect 635 21 643 25
rect 635 19 638 21
rect 640 19 643 21
rect 635 17 643 19
rect 645 24 652 26
rect 645 22 648 24
rect 650 22 652 24
rect 645 20 652 22
rect 645 17 650 20
<< pdif >>
rect 9 527 14 542
rect 7 525 14 527
rect 7 523 9 525
rect 11 523 14 525
rect 7 521 14 523
rect 9 515 14 521
rect 16 533 24 542
rect 16 531 19 533
rect 21 531 24 533
rect 16 524 24 531
rect 26 540 34 542
rect 26 538 29 540
rect 31 538 34 540
rect 26 533 34 538
rect 26 531 29 533
rect 31 531 34 533
rect 26 524 34 531
rect 36 526 50 542
rect 36 524 45 526
rect 47 524 50 526
rect 16 515 21 524
rect 38 519 50 524
rect 38 517 45 519
rect 47 517 50 519
rect 38 515 50 517
rect 52 540 59 542
rect 52 538 55 540
rect 57 538 59 540
rect 52 536 59 538
rect 52 515 57 536
rect 92 535 98 542
rect 71 526 78 535
rect 71 524 73 526
rect 75 524 78 526
rect 71 522 78 524
rect 80 533 88 535
rect 80 531 83 533
rect 85 531 88 533
rect 80 526 88 531
rect 80 524 83 526
rect 85 524 88 526
rect 80 522 88 524
rect 90 528 98 535
rect 90 526 93 528
rect 95 526 98 528
rect 90 524 98 526
rect 100 540 107 542
rect 100 538 103 540
rect 105 538 107 540
rect 100 533 107 538
rect 100 531 103 533
rect 105 531 107 533
rect 100 529 107 531
rect 100 524 105 529
rect 113 527 118 542
rect 111 525 118 527
rect 90 522 96 524
rect 111 523 113 525
rect 115 523 118 525
rect 111 521 118 523
rect 113 515 118 521
rect 120 533 128 542
rect 120 531 123 533
rect 125 531 128 533
rect 120 524 128 531
rect 130 540 138 542
rect 130 538 133 540
rect 135 538 138 540
rect 130 533 138 538
rect 130 531 133 533
rect 135 531 138 533
rect 130 524 138 531
rect 140 526 154 542
rect 140 524 149 526
rect 151 524 154 526
rect 120 515 125 524
rect 142 519 154 524
rect 142 517 149 519
rect 151 517 154 519
rect 142 515 154 517
rect 156 540 163 542
rect 156 538 159 540
rect 161 538 163 540
rect 156 536 163 538
rect 156 515 161 536
rect 196 535 202 542
rect 175 526 182 535
rect 175 524 177 526
rect 179 524 182 526
rect 175 522 182 524
rect 184 533 192 535
rect 184 531 187 533
rect 189 531 192 533
rect 184 526 192 531
rect 184 524 187 526
rect 189 524 192 526
rect 184 522 192 524
rect 194 528 202 535
rect 194 526 197 528
rect 199 526 202 528
rect 194 524 202 526
rect 204 540 211 542
rect 204 538 207 540
rect 209 538 211 540
rect 204 533 211 538
rect 234 536 242 543
rect 204 531 207 533
rect 209 531 211 533
rect 204 529 211 531
rect 204 524 209 529
rect 217 528 222 536
rect 215 526 222 528
rect 215 524 217 526
rect 219 524 222 526
rect 194 522 200 524
rect 215 522 222 524
rect 217 515 222 522
rect 224 515 229 536
rect 231 525 242 536
rect 244 538 249 543
rect 244 536 251 538
rect 244 534 247 536
rect 249 534 251 536
rect 244 529 251 534
rect 244 527 247 529
rect 249 527 251 529
rect 258 527 263 542
rect 244 525 251 527
rect 256 525 263 527
rect 231 519 240 525
rect 256 523 258 525
rect 260 523 263 525
rect 256 521 263 523
rect 231 517 236 519
rect 238 517 240 519
rect 231 515 240 517
rect 258 515 263 521
rect 265 533 273 542
rect 265 531 268 533
rect 270 531 273 533
rect 265 524 273 531
rect 275 540 283 542
rect 275 538 278 540
rect 280 538 283 540
rect 275 533 283 538
rect 275 531 278 533
rect 280 531 283 533
rect 275 524 283 531
rect 285 526 299 542
rect 285 524 294 526
rect 296 524 299 526
rect 265 515 270 524
rect 287 519 299 524
rect 287 517 294 519
rect 296 517 299 519
rect 287 515 299 517
rect 301 540 308 542
rect 301 538 304 540
rect 306 538 308 540
rect 301 536 308 538
rect 301 515 306 536
rect 341 535 347 542
rect 320 526 327 535
rect 320 524 322 526
rect 324 524 327 526
rect 320 522 327 524
rect 329 533 337 535
rect 329 531 332 533
rect 334 531 337 533
rect 329 526 337 531
rect 329 524 332 526
rect 334 524 337 526
rect 329 522 337 524
rect 339 528 347 535
rect 339 526 342 528
rect 344 526 347 528
rect 339 524 347 526
rect 349 540 356 542
rect 349 538 352 540
rect 354 538 356 540
rect 349 533 356 538
rect 379 536 387 543
rect 349 531 352 533
rect 354 531 356 533
rect 349 529 356 531
rect 349 524 354 529
rect 362 528 367 536
rect 360 526 367 528
rect 360 524 362 526
rect 364 524 367 526
rect 339 522 345 524
rect 360 522 367 524
rect 362 515 367 522
rect 369 515 374 536
rect 376 525 387 536
rect 389 538 394 543
rect 408 540 415 542
rect 408 538 410 540
rect 412 538 415 540
rect 389 536 396 538
rect 408 536 415 538
rect 389 534 392 536
rect 394 534 396 536
rect 389 529 396 534
rect 389 527 392 529
rect 394 527 396 529
rect 389 525 396 527
rect 376 519 385 525
rect 376 517 381 519
rect 383 517 385 519
rect 376 515 385 517
rect 410 515 415 536
rect 417 526 431 542
rect 417 524 420 526
rect 422 524 431 526
rect 433 540 441 542
rect 433 538 436 540
rect 438 538 441 540
rect 433 533 441 538
rect 433 531 436 533
rect 438 531 441 533
rect 433 524 441 531
rect 443 533 451 542
rect 443 531 446 533
rect 448 531 451 533
rect 443 524 451 531
rect 417 519 429 524
rect 417 517 420 519
rect 422 517 429 519
rect 417 515 429 517
rect 446 515 451 524
rect 453 527 458 542
rect 464 541 471 543
rect 464 539 466 541
rect 468 539 471 541
rect 464 537 471 539
rect 466 535 471 537
rect 473 535 479 543
rect 475 531 479 535
rect 528 541 535 543
rect 528 539 530 541
rect 532 539 535 541
rect 528 537 535 539
rect 530 535 535 537
rect 537 535 543 543
rect 510 531 515 533
rect 453 525 460 527
rect 475 527 481 531
rect 453 523 456 525
rect 458 523 460 525
rect 453 521 460 523
rect 453 515 458 521
rect 474 519 481 527
rect 474 517 476 519
rect 478 517 481 519
rect 474 515 481 517
rect 483 515 488 531
rect 490 529 498 531
rect 490 527 493 529
rect 495 527 498 529
rect 490 515 498 527
rect 500 515 505 531
rect 507 519 515 531
rect 507 517 510 519
rect 512 517 515 519
rect 507 515 515 517
rect 517 528 522 533
rect 539 531 543 535
rect 592 541 599 543
rect 592 539 594 541
rect 596 539 599 541
rect 592 537 599 539
rect 594 535 599 537
rect 601 535 607 543
rect 574 531 579 533
rect 517 526 524 528
rect 539 527 545 531
rect 517 524 520 526
rect 522 524 524 526
rect 517 522 524 524
rect 517 515 522 522
rect 538 519 545 527
rect 538 517 540 519
rect 542 517 545 519
rect 538 515 545 517
rect 547 515 552 531
rect 554 529 562 531
rect 554 527 557 529
rect 559 527 562 529
rect 554 515 562 527
rect 564 515 569 531
rect 571 519 579 531
rect 571 517 574 519
rect 576 517 579 519
rect 571 515 579 517
rect 581 528 586 533
rect 603 531 607 535
rect 638 531 643 533
rect 581 526 588 528
rect 603 527 609 531
rect 581 524 584 526
rect 586 524 588 526
rect 581 522 588 524
rect 581 515 586 522
rect 602 519 609 527
rect 602 517 604 519
rect 606 517 609 519
rect 602 515 609 517
rect 611 515 616 531
rect 618 529 626 531
rect 618 527 621 529
rect 623 527 626 529
rect 618 515 626 527
rect 628 515 633 531
rect 635 519 643 531
rect 635 517 638 519
rect 640 517 643 519
rect 635 515 643 517
rect 645 528 650 533
rect 645 526 652 528
rect 645 524 648 526
rect 650 524 652 526
rect 645 522 652 524
rect 645 515 650 522
rect 18 501 27 503
rect 18 499 20 501
rect 22 499 27 501
rect 18 493 27 499
rect 7 491 14 493
rect 7 489 9 491
rect 11 489 14 491
rect 7 484 14 489
rect 7 482 9 484
rect 11 482 14 484
rect 7 480 14 482
rect 9 475 14 480
rect 16 482 27 493
rect 29 482 34 503
rect 36 496 41 503
rect 36 494 43 496
rect 58 494 64 496
rect 36 492 39 494
rect 41 492 43 494
rect 36 490 43 492
rect 36 482 41 490
rect 49 489 54 494
rect 47 487 54 489
rect 47 485 49 487
rect 51 485 54 487
rect 16 475 24 482
rect 47 480 54 485
rect 47 478 49 480
rect 51 478 54 480
rect 47 476 54 478
rect 56 492 64 494
rect 56 490 59 492
rect 61 490 64 492
rect 56 483 64 490
rect 66 494 74 496
rect 66 492 69 494
rect 71 492 74 494
rect 66 487 74 492
rect 66 485 69 487
rect 71 485 74 487
rect 66 483 74 485
rect 76 494 83 496
rect 76 492 79 494
rect 81 492 83 494
rect 76 483 83 492
rect 56 476 62 483
rect 97 482 102 503
rect 95 480 102 482
rect 95 478 97 480
rect 99 478 102 480
rect 95 476 102 478
rect 104 501 116 503
rect 104 499 107 501
rect 109 499 116 501
rect 104 494 116 499
rect 133 494 138 503
rect 104 492 107 494
rect 109 492 118 494
rect 104 476 118 492
rect 120 487 128 494
rect 120 485 123 487
rect 125 485 128 487
rect 120 480 128 485
rect 120 478 123 480
rect 125 478 128 480
rect 120 476 128 478
rect 130 487 138 494
rect 130 485 133 487
rect 135 485 138 487
rect 130 476 138 485
rect 140 497 145 503
rect 140 495 147 497
rect 140 493 143 495
rect 145 493 147 495
rect 162 494 168 496
rect 140 491 147 493
rect 140 476 145 491
rect 153 489 158 494
rect 151 487 158 489
rect 151 485 153 487
rect 155 485 158 487
rect 151 480 158 485
rect 151 478 153 480
rect 155 478 158 480
rect 151 476 158 478
rect 160 492 168 494
rect 160 490 163 492
rect 165 490 168 492
rect 160 483 168 490
rect 170 494 178 496
rect 170 492 173 494
rect 175 492 178 494
rect 170 487 178 492
rect 170 485 173 487
rect 175 485 178 487
rect 170 483 178 485
rect 180 494 187 496
rect 180 492 183 494
rect 185 492 187 494
rect 180 483 187 492
rect 160 476 166 483
rect 201 482 206 503
rect 199 480 206 482
rect 199 478 201 480
rect 203 478 206 480
rect 199 476 206 478
rect 208 501 220 503
rect 208 499 211 501
rect 213 499 220 501
rect 208 494 220 499
rect 237 494 242 503
rect 208 492 211 494
rect 213 492 222 494
rect 208 476 222 492
rect 224 487 232 494
rect 224 485 227 487
rect 229 485 232 487
rect 224 480 232 485
rect 224 478 227 480
rect 229 478 232 480
rect 224 476 232 478
rect 234 487 242 494
rect 234 485 237 487
rect 239 485 242 487
rect 234 476 242 485
rect 244 497 249 503
rect 258 497 263 503
rect 244 495 251 497
rect 244 493 247 495
rect 249 493 251 495
rect 244 491 251 493
rect 256 495 263 497
rect 256 493 258 495
rect 260 493 263 495
rect 256 491 263 493
rect 244 476 249 491
rect 258 476 263 491
rect 265 494 270 503
rect 287 501 299 503
rect 287 499 294 501
rect 296 499 299 501
rect 287 494 299 499
rect 265 487 273 494
rect 265 485 268 487
rect 270 485 273 487
rect 265 476 273 485
rect 275 487 283 494
rect 275 485 278 487
rect 280 485 283 487
rect 275 480 283 485
rect 275 478 278 480
rect 280 478 283 480
rect 275 476 283 478
rect 285 492 294 494
rect 296 492 299 494
rect 285 476 299 492
rect 301 482 306 503
rect 320 494 327 496
rect 320 492 322 494
rect 324 492 327 494
rect 320 483 327 492
rect 329 494 337 496
rect 329 492 332 494
rect 334 492 337 494
rect 329 487 337 492
rect 329 485 332 487
rect 334 485 337 487
rect 329 483 337 485
rect 339 494 345 496
rect 362 496 367 503
rect 360 494 367 496
rect 339 492 347 494
rect 339 490 342 492
rect 344 490 347 492
rect 339 483 347 490
rect 301 480 308 482
rect 301 478 304 480
rect 306 478 308 480
rect 301 476 308 478
rect 341 476 347 483
rect 349 489 354 494
rect 360 492 362 494
rect 364 492 367 494
rect 360 490 367 492
rect 349 487 356 489
rect 349 485 352 487
rect 354 485 356 487
rect 349 480 356 485
rect 362 482 367 490
rect 369 482 374 503
rect 376 501 385 503
rect 376 499 381 501
rect 383 499 385 501
rect 376 493 385 499
rect 376 482 387 493
rect 349 478 352 480
rect 354 478 356 480
rect 349 476 356 478
rect 379 475 387 482
rect 389 491 396 493
rect 389 489 392 491
rect 394 489 396 491
rect 389 484 396 489
rect 389 482 392 484
rect 394 482 396 484
rect 410 482 415 503
rect 389 480 396 482
rect 408 480 415 482
rect 389 475 394 480
rect 408 478 410 480
rect 412 478 415 480
rect 408 476 415 478
rect 417 501 429 503
rect 417 499 420 501
rect 422 499 429 501
rect 417 494 429 499
rect 446 494 451 503
rect 417 492 420 494
rect 422 492 431 494
rect 417 476 431 492
rect 433 487 441 494
rect 433 485 436 487
rect 438 485 441 487
rect 433 480 441 485
rect 433 478 436 480
rect 438 478 441 480
rect 433 476 441 478
rect 443 487 451 494
rect 443 485 446 487
rect 448 485 451 487
rect 443 476 451 485
rect 453 497 458 503
rect 474 501 481 503
rect 474 499 476 501
rect 478 499 481 501
rect 453 495 460 497
rect 453 493 456 495
rect 458 493 460 495
rect 453 491 460 493
rect 453 476 458 491
rect 474 491 481 499
rect 475 487 481 491
rect 483 487 488 503
rect 490 491 498 503
rect 490 489 493 491
rect 495 489 498 491
rect 490 487 498 489
rect 500 487 505 503
rect 507 501 515 503
rect 507 499 510 501
rect 512 499 515 501
rect 507 487 515 499
rect 475 483 479 487
rect 466 481 471 483
rect 464 479 471 481
rect 464 477 466 479
rect 468 477 471 479
rect 464 475 471 477
rect 473 475 479 483
rect 510 485 515 487
rect 517 496 522 503
rect 538 501 545 503
rect 538 499 540 501
rect 542 499 545 501
rect 517 494 524 496
rect 517 492 520 494
rect 522 492 524 494
rect 517 490 524 492
rect 538 491 545 499
rect 517 485 522 490
rect 539 487 545 491
rect 547 487 552 503
rect 554 491 562 503
rect 554 489 557 491
rect 559 489 562 491
rect 554 487 562 489
rect 564 487 569 503
rect 571 501 579 503
rect 571 499 574 501
rect 576 499 579 501
rect 571 487 579 499
rect 539 483 543 487
rect 530 481 535 483
rect 528 479 535 481
rect 528 477 530 479
rect 532 477 535 479
rect 528 475 535 477
rect 537 475 543 483
rect 574 485 579 487
rect 581 496 586 503
rect 602 501 609 503
rect 602 499 604 501
rect 606 499 609 501
rect 581 494 588 496
rect 581 492 584 494
rect 586 492 588 494
rect 581 490 588 492
rect 602 491 609 499
rect 581 485 586 490
rect 603 487 609 491
rect 611 487 616 503
rect 618 491 626 503
rect 618 489 621 491
rect 623 489 626 491
rect 618 487 626 489
rect 628 487 633 503
rect 635 501 643 503
rect 635 499 638 501
rect 640 499 643 501
rect 635 487 643 499
rect 603 483 607 487
rect 594 481 599 483
rect 592 479 599 481
rect 592 477 594 479
rect 596 477 599 479
rect 592 475 599 477
rect 601 475 607 483
rect 638 485 643 487
rect 645 496 650 503
rect 645 494 652 496
rect 645 492 648 494
rect 650 492 652 494
rect 645 490 652 492
rect 645 485 650 490
rect 9 383 14 398
rect 7 381 14 383
rect 7 379 9 381
rect 11 379 14 381
rect 7 377 14 379
rect 9 371 14 377
rect 16 389 24 398
rect 16 387 19 389
rect 21 387 24 389
rect 16 380 24 387
rect 26 396 34 398
rect 26 394 29 396
rect 31 394 34 396
rect 26 389 34 394
rect 26 387 29 389
rect 31 387 34 389
rect 26 380 34 387
rect 36 382 50 398
rect 36 380 45 382
rect 47 380 50 382
rect 16 371 21 380
rect 38 375 50 380
rect 38 373 45 375
rect 47 373 50 375
rect 38 371 50 373
rect 52 396 59 398
rect 52 394 55 396
rect 57 394 59 396
rect 52 392 59 394
rect 52 371 57 392
rect 92 391 98 398
rect 71 382 78 391
rect 71 380 73 382
rect 75 380 78 382
rect 71 378 78 380
rect 80 389 88 391
rect 80 387 83 389
rect 85 387 88 389
rect 80 382 88 387
rect 80 380 83 382
rect 85 380 88 382
rect 80 378 88 380
rect 90 384 98 391
rect 90 382 93 384
rect 95 382 98 384
rect 90 380 98 382
rect 100 396 107 398
rect 100 394 103 396
rect 105 394 107 396
rect 100 389 107 394
rect 100 387 103 389
rect 105 387 107 389
rect 100 385 107 387
rect 100 380 105 385
rect 113 383 118 398
rect 111 381 118 383
rect 90 378 96 380
rect 111 379 113 381
rect 115 379 118 381
rect 111 377 118 379
rect 113 371 118 377
rect 120 389 128 398
rect 120 387 123 389
rect 125 387 128 389
rect 120 380 128 387
rect 130 396 138 398
rect 130 394 133 396
rect 135 394 138 396
rect 130 389 138 394
rect 130 387 133 389
rect 135 387 138 389
rect 130 380 138 387
rect 140 382 154 398
rect 140 380 149 382
rect 151 380 154 382
rect 120 371 125 380
rect 142 375 154 380
rect 142 373 149 375
rect 151 373 154 375
rect 142 371 154 373
rect 156 396 163 398
rect 156 394 159 396
rect 161 394 163 396
rect 156 392 163 394
rect 156 371 161 392
rect 196 391 202 398
rect 175 382 182 391
rect 175 380 177 382
rect 179 380 182 382
rect 175 378 182 380
rect 184 389 192 391
rect 184 387 187 389
rect 189 387 192 389
rect 184 382 192 387
rect 184 380 187 382
rect 189 380 192 382
rect 184 378 192 380
rect 194 384 202 391
rect 194 382 197 384
rect 199 382 202 384
rect 194 380 202 382
rect 204 396 211 398
rect 204 394 207 396
rect 209 394 211 396
rect 204 389 211 394
rect 234 392 242 399
rect 204 387 207 389
rect 209 387 211 389
rect 204 385 211 387
rect 204 380 209 385
rect 217 384 222 392
rect 215 382 222 384
rect 215 380 217 382
rect 219 380 222 382
rect 194 378 200 380
rect 215 378 222 380
rect 217 371 222 378
rect 224 371 229 392
rect 231 381 242 392
rect 244 394 249 399
rect 244 392 251 394
rect 244 390 247 392
rect 249 390 251 392
rect 244 385 251 390
rect 244 383 247 385
rect 249 383 251 385
rect 258 383 263 398
rect 244 381 251 383
rect 256 381 263 383
rect 231 375 240 381
rect 256 379 258 381
rect 260 379 263 381
rect 256 377 263 379
rect 231 373 236 375
rect 238 373 240 375
rect 231 371 240 373
rect 258 371 263 377
rect 265 389 273 398
rect 265 387 268 389
rect 270 387 273 389
rect 265 380 273 387
rect 275 396 283 398
rect 275 394 278 396
rect 280 394 283 396
rect 275 389 283 394
rect 275 387 278 389
rect 280 387 283 389
rect 275 380 283 387
rect 285 382 299 398
rect 285 380 294 382
rect 296 380 299 382
rect 265 371 270 380
rect 287 375 299 380
rect 287 373 294 375
rect 296 373 299 375
rect 287 371 299 373
rect 301 396 308 398
rect 301 394 304 396
rect 306 394 308 396
rect 301 392 308 394
rect 301 371 306 392
rect 341 391 347 398
rect 320 382 327 391
rect 320 380 322 382
rect 324 380 327 382
rect 320 378 327 380
rect 329 389 337 391
rect 329 387 332 389
rect 334 387 337 389
rect 329 382 337 387
rect 329 380 332 382
rect 334 380 337 382
rect 329 378 337 380
rect 339 384 347 391
rect 339 382 342 384
rect 344 382 347 384
rect 339 380 347 382
rect 349 396 356 398
rect 349 394 352 396
rect 354 394 356 396
rect 349 389 356 394
rect 379 392 387 399
rect 349 387 352 389
rect 354 387 356 389
rect 349 385 356 387
rect 349 380 354 385
rect 362 384 367 392
rect 360 382 367 384
rect 360 380 362 382
rect 364 380 367 382
rect 339 378 345 380
rect 360 378 367 380
rect 362 371 367 378
rect 369 371 374 392
rect 376 381 387 392
rect 389 394 394 399
rect 408 396 415 398
rect 408 394 410 396
rect 412 394 415 396
rect 389 392 396 394
rect 408 392 415 394
rect 389 390 392 392
rect 394 390 396 392
rect 389 385 396 390
rect 389 383 392 385
rect 394 383 396 385
rect 389 381 396 383
rect 376 375 385 381
rect 376 373 381 375
rect 383 373 385 375
rect 376 371 385 373
rect 410 371 415 392
rect 417 382 431 398
rect 417 380 420 382
rect 422 380 431 382
rect 433 396 441 398
rect 433 394 436 396
rect 438 394 441 396
rect 433 389 441 394
rect 433 387 436 389
rect 438 387 441 389
rect 433 380 441 387
rect 443 389 451 398
rect 443 387 446 389
rect 448 387 451 389
rect 443 380 451 387
rect 417 375 429 380
rect 417 373 420 375
rect 422 373 429 375
rect 417 371 429 373
rect 446 371 451 380
rect 453 383 458 398
rect 464 397 471 399
rect 464 395 466 397
rect 468 395 471 397
rect 464 393 471 395
rect 466 391 471 393
rect 473 391 479 399
rect 475 387 479 391
rect 528 397 535 399
rect 528 395 530 397
rect 532 395 535 397
rect 528 393 535 395
rect 530 391 535 393
rect 537 391 543 399
rect 510 387 515 389
rect 453 381 460 383
rect 475 383 481 387
rect 453 379 456 381
rect 458 379 460 381
rect 453 377 460 379
rect 453 371 458 377
rect 474 375 481 383
rect 474 373 476 375
rect 478 373 481 375
rect 474 371 481 373
rect 483 371 488 387
rect 490 385 498 387
rect 490 383 493 385
rect 495 383 498 385
rect 490 371 498 383
rect 500 371 505 387
rect 507 375 515 387
rect 507 373 510 375
rect 512 373 515 375
rect 507 371 515 373
rect 517 384 522 389
rect 539 387 543 391
rect 592 397 599 399
rect 592 395 594 397
rect 596 395 599 397
rect 592 393 599 395
rect 594 391 599 393
rect 601 391 607 399
rect 574 387 579 389
rect 517 382 524 384
rect 539 383 545 387
rect 517 380 520 382
rect 522 380 524 382
rect 517 378 524 380
rect 517 371 522 378
rect 538 375 545 383
rect 538 373 540 375
rect 542 373 545 375
rect 538 371 545 373
rect 547 371 552 387
rect 554 385 562 387
rect 554 383 557 385
rect 559 383 562 385
rect 554 371 562 383
rect 564 371 569 387
rect 571 375 579 387
rect 571 373 574 375
rect 576 373 579 375
rect 571 371 579 373
rect 581 384 586 389
rect 603 387 607 391
rect 638 387 643 389
rect 581 382 588 384
rect 603 383 609 387
rect 581 380 584 382
rect 586 380 588 382
rect 581 378 588 380
rect 581 371 586 378
rect 602 375 609 383
rect 602 373 604 375
rect 606 373 609 375
rect 602 371 609 373
rect 611 371 616 387
rect 618 385 626 387
rect 618 383 621 385
rect 623 383 626 385
rect 618 371 626 383
rect 628 371 633 387
rect 635 375 643 387
rect 635 373 638 375
rect 640 373 643 375
rect 635 371 643 373
rect 645 384 650 389
rect 645 382 652 384
rect 645 380 648 382
rect 650 380 652 382
rect 645 378 652 380
rect 645 371 650 378
rect 18 357 27 359
rect 18 355 20 357
rect 22 355 27 357
rect 18 349 27 355
rect 7 347 14 349
rect 7 345 9 347
rect 11 345 14 347
rect 7 340 14 345
rect 7 338 9 340
rect 11 338 14 340
rect 7 336 14 338
rect 9 331 14 336
rect 16 338 27 349
rect 29 338 34 359
rect 36 352 41 359
rect 36 350 43 352
rect 58 350 64 352
rect 36 348 39 350
rect 41 348 43 350
rect 36 346 43 348
rect 36 338 41 346
rect 49 345 54 350
rect 47 343 54 345
rect 47 341 49 343
rect 51 341 54 343
rect 16 331 24 338
rect 47 336 54 341
rect 47 334 49 336
rect 51 334 54 336
rect 47 332 54 334
rect 56 348 64 350
rect 56 346 59 348
rect 61 346 64 348
rect 56 339 64 346
rect 66 350 74 352
rect 66 348 69 350
rect 71 348 74 350
rect 66 343 74 348
rect 66 341 69 343
rect 71 341 74 343
rect 66 339 74 341
rect 76 350 83 352
rect 76 348 79 350
rect 81 348 83 350
rect 76 339 83 348
rect 56 332 62 339
rect 97 338 102 359
rect 95 336 102 338
rect 95 334 97 336
rect 99 334 102 336
rect 95 332 102 334
rect 104 357 116 359
rect 104 355 107 357
rect 109 355 116 357
rect 104 350 116 355
rect 133 350 138 359
rect 104 348 107 350
rect 109 348 118 350
rect 104 332 118 348
rect 120 343 128 350
rect 120 341 123 343
rect 125 341 128 343
rect 120 336 128 341
rect 120 334 123 336
rect 125 334 128 336
rect 120 332 128 334
rect 130 343 138 350
rect 130 341 133 343
rect 135 341 138 343
rect 130 332 138 341
rect 140 353 145 359
rect 140 351 147 353
rect 140 349 143 351
rect 145 349 147 351
rect 162 350 168 352
rect 140 347 147 349
rect 140 332 145 347
rect 153 345 158 350
rect 151 343 158 345
rect 151 341 153 343
rect 155 341 158 343
rect 151 336 158 341
rect 151 334 153 336
rect 155 334 158 336
rect 151 332 158 334
rect 160 348 168 350
rect 160 346 163 348
rect 165 346 168 348
rect 160 339 168 346
rect 170 350 178 352
rect 170 348 173 350
rect 175 348 178 350
rect 170 343 178 348
rect 170 341 173 343
rect 175 341 178 343
rect 170 339 178 341
rect 180 350 187 352
rect 180 348 183 350
rect 185 348 187 350
rect 180 339 187 348
rect 160 332 166 339
rect 201 338 206 359
rect 199 336 206 338
rect 199 334 201 336
rect 203 334 206 336
rect 199 332 206 334
rect 208 357 220 359
rect 208 355 211 357
rect 213 355 220 357
rect 208 350 220 355
rect 237 350 242 359
rect 208 348 211 350
rect 213 348 222 350
rect 208 332 222 348
rect 224 343 232 350
rect 224 341 227 343
rect 229 341 232 343
rect 224 336 232 341
rect 224 334 227 336
rect 229 334 232 336
rect 224 332 232 334
rect 234 343 242 350
rect 234 341 237 343
rect 239 341 242 343
rect 234 332 242 341
rect 244 353 249 359
rect 258 353 263 359
rect 244 351 251 353
rect 244 349 247 351
rect 249 349 251 351
rect 244 347 251 349
rect 256 351 263 353
rect 256 349 258 351
rect 260 349 263 351
rect 256 347 263 349
rect 244 332 249 347
rect 258 332 263 347
rect 265 350 270 359
rect 287 357 299 359
rect 287 355 294 357
rect 296 355 299 357
rect 287 350 299 355
rect 265 343 273 350
rect 265 341 268 343
rect 270 341 273 343
rect 265 332 273 341
rect 275 343 283 350
rect 275 341 278 343
rect 280 341 283 343
rect 275 336 283 341
rect 275 334 278 336
rect 280 334 283 336
rect 275 332 283 334
rect 285 348 294 350
rect 296 348 299 350
rect 285 332 299 348
rect 301 338 306 359
rect 320 350 327 352
rect 320 348 322 350
rect 324 348 327 350
rect 320 339 327 348
rect 329 350 337 352
rect 329 348 332 350
rect 334 348 337 350
rect 329 343 337 348
rect 329 341 332 343
rect 334 341 337 343
rect 329 339 337 341
rect 339 350 345 352
rect 362 352 367 359
rect 360 350 367 352
rect 339 348 347 350
rect 339 346 342 348
rect 344 346 347 348
rect 339 339 347 346
rect 301 336 308 338
rect 301 334 304 336
rect 306 334 308 336
rect 301 332 308 334
rect 341 332 347 339
rect 349 345 354 350
rect 360 348 362 350
rect 364 348 367 350
rect 360 346 367 348
rect 349 343 356 345
rect 349 341 352 343
rect 354 341 356 343
rect 349 336 356 341
rect 362 338 367 346
rect 369 338 374 359
rect 376 357 385 359
rect 376 355 381 357
rect 383 355 385 357
rect 376 349 385 355
rect 376 338 387 349
rect 349 334 352 336
rect 354 334 356 336
rect 349 332 356 334
rect 379 331 387 338
rect 389 347 396 349
rect 389 345 392 347
rect 394 345 396 347
rect 389 340 396 345
rect 389 338 392 340
rect 394 338 396 340
rect 410 338 415 359
rect 389 336 396 338
rect 408 336 415 338
rect 389 331 394 336
rect 408 334 410 336
rect 412 334 415 336
rect 408 332 415 334
rect 417 357 429 359
rect 417 355 420 357
rect 422 355 429 357
rect 417 350 429 355
rect 446 350 451 359
rect 417 348 420 350
rect 422 348 431 350
rect 417 332 431 348
rect 433 343 441 350
rect 433 341 436 343
rect 438 341 441 343
rect 433 336 441 341
rect 433 334 436 336
rect 438 334 441 336
rect 433 332 441 334
rect 443 343 451 350
rect 443 341 446 343
rect 448 341 451 343
rect 443 332 451 341
rect 453 353 458 359
rect 474 357 481 359
rect 474 355 476 357
rect 478 355 481 357
rect 453 351 460 353
rect 453 349 456 351
rect 458 349 460 351
rect 453 347 460 349
rect 453 332 458 347
rect 474 347 481 355
rect 475 343 481 347
rect 483 343 488 359
rect 490 347 498 359
rect 490 345 493 347
rect 495 345 498 347
rect 490 343 498 345
rect 500 343 505 359
rect 507 357 515 359
rect 507 355 510 357
rect 512 355 515 357
rect 507 343 515 355
rect 475 339 479 343
rect 466 337 471 339
rect 464 335 471 337
rect 464 333 466 335
rect 468 333 471 335
rect 464 331 471 333
rect 473 331 479 339
rect 510 341 515 343
rect 517 352 522 359
rect 538 357 545 359
rect 538 355 540 357
rect 542 355 545 357
rect 517 350 524 352
rect 517 348 520 350
rect 522 348 524 350
rect 517 346 524 348
rect 538 347 545 355
rect 517 341 522 346
rect 539 343 545 347
rect 547 343 552 359
rect 554 347 562 359
rect 554 345 557 347
rect 559 345 562 347
rect 554 343 562 345
rect 564 343 569 359
rect 571 357 579 359
rect 571 355 574 357
rect 576 355 579 357
rect 571 343 579 355
rect 539 339 543 343
rect 530 337 535 339
rect 528 335 535 337
rect 528 333 530 335
rect 532 333 535 335
rect 528 331 535 333
rect 537 331 543 339
rect 574 341 579 343
rect 581 352 586 359
rect 602 357 609 359
rect 602 355 604 357
rect 606 355 609 357
rect 581 350 588 352
rect 581 348 584 350
rect 586 348 588 350
rect 581 346 588 348
rect 602 347 609 355
rect 581 341 586 346
rect 603 343 609 347
rect 611 343 616 359
rect 618 347 626 359
rect 618 345 621 347
rect 623 345 626 347
rect 618 343 626 345
rect 628 343 633 359
rect 635 357 643 359
rect 635 355 638 357
rect 640 355 643 357
rect 635 343 643 355
rect 603 339 607 343
rect 594 337 599 339
rect 592 335 599 337
rect 592 333 594 335
rect 596 333 599 335
rect 592 331 599 333
rect 601 331 607 339
rect 638 341 643 343
rect 645 352 650 359
rect 645 350 652 352
rect 645 348 648 350
rect 650 348 652 350
rect 645 346 652 348
rect 645 341 650 346
rect 9 239 14 254
rect 7 237 14 239
rect 7 235 9 237
rect 11 235 14 237
rect 7 233 14 235
rect 9 227 14 233
rect 16 245 24 254
rect 16 243 19 245
rect 21 243 24 245
rect 16 236 24 243
rect 26 252 34 254
rect 26 250 29 252
rect 31 250 34 252
rect 26 245 34 250
rect 26 243 29 245
rect 31 243 34 245
rect 26 236 34 243
rect 36 238 50 254
rect 36 236 45 238
rect 47 236 50 238
rect 16 227 21 236
rect 38 231 50 236
rect 38 229 45 231
rect 47 229 50 231
rect 38 227 50 229
rect 52 252 59 254
rect 52 250 55 252
rect 57 250 59 252
rect 52 248 59 250
rect 52 227 57 248
rect 92 247 98 254
rect 71 238 78 247
rect 71 236 73 238
rect 75 236 78 238
rect 71 234 78 236
rect 80 245 88 247
rect 80 243 83 245
rect 85 243 88 245
rect 80 238 88 243
rect 80 236 83 238
rect 85 236 88 238
rect 80 234 88 236
rect 90 240 98 247
rect 90 238 93 240
rect 95 238 98 240
rect 90 236 98 238
rect 100 252 107 254
rect 100 250 103 252
rect 105 250 107 252
rect 100 245 107 250
rect 100 243 103 245
rect 105 243 107 245
rect 100 241 107 243
rect 100 236 105 241
rect 113 239 118 254
rect 111 237 118 239
rect 90 234 96 236
rect 111 235 113 237
rect 115 235 118 237
rect 111 233 118 235
rect 113 227 118 233
rect 120 245 128 254
rect 120 243 123 245
rect 125 243 128 245
rect 120 236 128 243
rect 130 252 138 254
rect 130 250 133 252
rect 135 250 138 252
rect 130 245 138 250
rect 130 243 133 245
rect 135 243 138 245
rect 130 236 138 243
rect 140 238 154 254
rect 140 236 149 238
rect 151 236 154 238
rect 120 227 125 236
rect 142 231 154 236
rect 142 229 149 231
rect 151 229 154 231
rect 142 227 154 229
rect 156 252 163 254
rect 156 250 159 252
rect 161 250 163 252
rect 156 248 163 250
rect 156 227 161 248
rect 196 247 202 254
rect 175 238 182 247
rect 175 236 177 238
rect 179 236 182 238
rect 175 234 182 236
rect 184 245 192 247
rect 184 243 187 245
rect 189 243 192 245
rect 184 238 192 243
rect 184 236 187 238
rect 189 236 192 238
rect 184 234 192 236
rect 194 240 202 247
rect 194 238 197 240
rect 199 238 202 240
rect 194 236 202 238
rect 204 252 211 254
rect 204 250 207 252
rect 209 250 211 252
rect 204 245 211 250
rect 234 248 242 255
rect 204 243 207 245
rect 209 243 211 245
rect 204 241 211 243
rect 204 236 209 241
rect 217 240 222 248
rect 215 238 222 240
rect 215 236 217 238
rect 219 236 222 238
rect 194 234 200 236
rect 215 234 222 236
rect 217 227 222 234
rect 224 227 229 248
rect 231 237 242 248
rect 244 250 249 255
rect 244 248 251 250
rect 244 246 247 248
rect 249 246 251 248
rect 244 241 251 246
rect 244 239 247 241
rect 249 239 251 241
rect 258 239 263 254
rect 244 237 251 239
rect 256 237 263 239
rect 231 231 240 237
rect 256 235 258 237
rect 260 235 263 237
rect 256 233 263 235
rect 231 229 236 231
rect 238 229 240 231
rect 231 227 240 229
rect 258 227 263 233
rect 265 245 273 254
rect 265 243 268 245
rect 270 243 273 245
rect 265 236 273 243
rect 275 252 283 254
rect 275 250 278 252
rect 280 250 283 252
rect 275 245 283 250
rect 275 243 278 245
rect 280 243 283 245
rect 275 236 283 243
rect 285 238 299 254
rect 285 236 294 238
rect 296 236 299 238
rect 265 227 270 236
rect 287 231 299 236
rect 287 229 294 231
rect 296 229 299 231
rect 287 227 299 229
rect 301 252 308 254
rect 301 250 304 252
rect 306 250 308 252
rect 301 248 308 250
rect 301 227 306 248
rect 341 247 347 254
rect 320 238 327 247
rect 320 236 322 238
rect 324 236 327 238
rect 320 234 327 236
rect 329 245 337 247
rect 329 243 332 245
rect 334 243 337 245
rect 329 238 337 243
rect 329 236 332 238
rect 334 236 337 238
rect 329 234 337 236
rect 339 240 347 247
rect 339 238 342 240
rect 344 238 347 240
rect 339 236 347 238
rect 349 252 356 254
rect 349 250 352 252
rect 354 250 356 252
rect 349 245 356 250
rect 379 248 387 255
rect 349 243 352 245
rect 354 243 356 245
rect 349 241 356 243
rect 349 236 354 241
rect 362 240 367 248
rect 360 238 367 240
rect 360 236 362 238
rect 364 236 367 238
rect 339 234 345 236
rect 360 234 367 236
rect 362 227 367 234
rect 369 227 374 248
rect 376 237 387 248
rect 389 250 394 255
rect 408 252 415 254
rect 408 250 410 252
rect 412 250 415 252
rect 389 248 396 250
rect 408 248 415 250
rect 389 246 392 248
rect 394 246 396 248
rect 389 241 396 246
rect 389 239 392 241
rect 394 239 396 241
rect 389 237 396 239
rect 376 231 385 237
rect 376 229 381 231
rect 383 229 385 231
rect 376 227 385 229
rect 410 227 415 248
rect 417 238 431 254
rect 417 236 420 238
rect 422 236 431 238
rect 433 252 441 254
rect 433 250 436 252
rect 438 250 441 252
rect 433 245 441 250
rect 433 243 436 245
rect 438 243 441 245
rect 433 236 441 243
rect 443 245 451 254
rect 443 243 446 245
rect 448 243 451 245
rect 443 236 451 243
rect 417 231 429 236
rect 417 229 420 231
rect 422 229 429 231
rect 417 227 429 229
rect 446 227 451 236
rect 453 239 458 254
rect 464 253 471 255
rect 464 251 466 253
rect 468 251 471 253
rect 464 249 471 251
rect 466 247 471 249
rect 473 247 479 255
rect 475 243 479 247
rect 528 253 535 255
rect 528 251 530 253
rect 532 251 535 253
rect 528 249 535 251
rect 530 247 535 249
rect 537 247 543 255
rect 510 243 515 245
rect 453 237 460 239
rect 475 239 481 243
rect 453 235 456 237
rect 458 235 460 237
rect 453 233 460 235
rect 453 227 458 233
rect 474 231 481 239
rect 474 229 476 231
rect 478 229 481 231
rect 474 227 481 229
rect 483 227 488 243
rect 490 241 498 243
rect 490 239 493 241
rect 495 239 498 241
rect 490 227 498 239
rect 500 227 505 243
rect 507 231 515 243
rect 507 229 510 231
rect 512 229 515 231
rect 507 227 515 229
rect 517 240 522 245
rect 539 243 543 247
rect 592 253 599 255
rect 592 251 594 253
rect 596 251 599 253
rect 592 249 599 251
rect 594 247 599 249
rect 601 247 607 255
rect 574 243 579 245
rect 517 238 524 240
rect 539 239 545 243
rect 517 236 520 238
rect 522 236 524 238
rect 517 234 524 236
rect 517 227 522 234
rect 538 231 545 239
rect 538 229 540 231
rect 542 229 545 231
rect 538 227 545 229
rect 547 227 552 243
rect 554 241 562 243
rect 554 239 557 241
rect 559 239 562 241
rect 554 227 562 239
rect 564 227 569 243
rect 571 231 579 243
rect 571 229 574 231
rect 576 229 579 231
rect 571 227 579 229
rect 581 240 586 245
rect 603 243 607 247
rect 638 243 643 245
rect 581 238 588 240
rect 603 239 609 243
rect 581 236 584 238
rect 586 236 588 238
rect 581 234 588 236
rect 581 227 586 234
rect 602 231 609 239
rect 602 229 604 231
rect 606 229 609 231
rect 602 227 609 229
rect 611 227 616 243
rect 618 241 626 243
rect 618 239 621 241
rect 623 239 626 241
rect 618 227 626 239
rect 628 227 633 243
rect 635 231 643 243
rect 635 229 638 231
rect 640 229 643 231
rect 635 227 643 229
rect 645 240 650 245
rect 645 238 652 240
rect 645 236 648 238
rect 650 236 652 238
rect 645 234 652 236
rect 645 227 650 234
rect 18 213 27 215
rect 18 211 20 213
rect 22 211 27 213
rect 18 205 27 211
rect 7 203 14 205
rect 7 201 9 203
rect 11 201 14 203
rect 7 196 14 201
rect 7 194 9 196
rect 11 194 14 196
rect 7 192 14 194
rect 9 187 14 192
rect 16 194 27 205
rect 29 194 34 215
rect 36 208 41 215
rect 36 206 43 208
rect 58 206 64 208
rect 36 204 39 206
rect 41 204 43 206
rect 36 202 43 204
rect 36 194 41 202
rect 49 201 54 206
rect 47 199 54 201
rect 47 197 49 199
rect 51 197 54 199
rect 16 187 24 194
rect 47 192 54 197
rect 47 190 49 192
rect 51 190 54 192
rect 47 188 54 190
rect 56 204 64 206
rect 56 202 59 204
rect 61 202 64 204
rect 56 195 64 202
rect 66 206 74 208
rect 66 204 69 206
rect 71 204 74 206
rect 66 199 74 204
rect 66 197 69 199
rect 71 197 74 199
rect 66 195 74 197
rect 76 206 83 208
rect 76 204 79 206
rect 81 204 83 206
rect 76 195 83 204
rect 56 188 62 195
rect 97 194 102 215
rect 95 192 102 194
rect 95 190 97 192
rect 99 190 102 192
rect 95 188 102 190
rect 104 213 116 215
rect 104 211 107 213
rect 109 211 116 213
rect 104 206 116 211
rect 133 206 138 215
rect 104 204 107 206
rect 109 204 118 206
rect 104 188 118 204
rect 120 199 128 206
rect 120 197 123 199
rect 125 197 128 199
rect 120 192 128 197
rect 120 190 123 192
rect 125 190 128 192
rect 120 188 128 190
rect 130 199 138 206
rect 130 197 133 199
rect 135 197 138 199
rect 130 188 138 197
rect 140 209 145 215
rect 140 207 147 209
rect 140 205 143 207
rect 145 205 147 207
rect 162 206 168 208
rect 140 203 147 205
rect 140 188 145 203
rect 153 201 158 206
rect 151 199 158 201
rect 151 197 153 199
rect 155 197 158 199
rect 151 192 158 197
rect 151 190 153 192
rect 155 190 158 192
rect 151 188 158 190
rect 160 204 168 206
rect 160 202 163 204
rect 165 202 168 204
rect 160 195 168 202
rect 170 206 178 208
rect 170 204 173 206
rect 175 204 178 206
rect 170 199 178 204
rect 170 197 173 199
rect 175 197 178 199
rect 170 195 178 197
rect 180 206 187 208
rect 180 204 183 206
rect 185 204 187 206
rect 180 195 187 204
rect 160 188 166 195
rect 201 194 206 215
rect 199 192 206 194
rect 199 190 201 192
rect 203 190 206 192
rect 199 188 206 190
rect 208 213 220 215
rect 208 211 211 213
rect 213 211 220 213
rect 208 206 220 211
rect 237 206 242 215
rect 208 204 211 206
rect 213 204 222 206
rect 208 188 222 204
rect 224 199 232 206
rect 224 197 227 199
rect 229 197 232 199
rect 224 192 232 197
rect 224 190 227 192
rect 229 190 232 192
rect 224 188 232 190
rect 234 199 242 206
rect 234 197 237 199
rect 239 197 242 199
rect 234 188 242 197
rect 244 209 249 215
rect 258 209 263 215
rect 244 207 251 209
rect 244 205 247 207
rect 249 205 251 207
rect 244 203 251 205
rect 256 207 263 209
rect 256 205 258 207
rect 260 205 263 207
rect 256 203 263 205
rect 244 188 249 203
rect 258 188 263 203
rect 265 206 270 215
rect 287 213 299 215
rect 287 211 294 213
rect 296 211 299 213
rect 287 206 299 211
rect 265 199 273 206
rect 265 197 268 199
rect 270 197 273 199
rect 265 188 273 197
rect 275 199 283 206
rect 275 197 278 199
rect 280 197 283 199
rect 275 192 283 197
rect 275 190 278 192
rect 280 190 283 192
rect 275 188 283 190
rect 285 204 294 206
rect 296 204 299 206
rect 285 188 299 204
rect 301 194 306 215
rect 320 206 327 208
rect 320 204 322 206
rect 324 204 327 206
rect 320 195 327 204
rect 329 206 337 208
rect 329 204 332 206
rect 334 204 337 206
rect 329 199 337 204
rect 329 197 332 199
rect 334 197 337 199
rect 329 195 337 197
rect 339 206 345 208
rect 362 208 367 215
rect 360 206 367 208
rect 339 204 347 206
rect 339 202 342 204
rect 344 202 347 204
rect 339 195 347 202
rect 301 192 308 194
rect 301 190 304 192
rect 306 190 308 192
rect 301 188 308 190
rect 341 188 347 195
rect 349 201 354 206
rect 360 204 362 206
rect 364 204 367 206
rect 360 202 367 204
rect 349 199 356 201
rect 349 197 352 199
rect 354 197 356 199
rect 349 192 356 197
rect 362 194 367 202
rect 369 194 374 215
rect 376 213 385 215
rect 376 211 381 213
rect 383 211 385 213
rect 376 205 385 211
rect 376 194 387 205
rect 349 190 352 192
rect 354 190 356 192
rect 349 188 356 190
rect 379 187 387 194
rect 389 203 396 205
rect 389 201 392 203
rect 394 201 396 203
rect 389 196 396 201
rect 389 194 392 196
rect 394 194 396 196
rect 410 194 415 215
rect 389 192 396 194
rect 408 192 415 194
rect 389 187 394 192
rect 408 190 410 192
rect 412 190 415 192
rect 408 188 415 190
rect 417 213 429 215
rect 417 211 420 213
rect 422 211 429 213
rect 417 206 429 211
rect 446 206 451 215
rect 417 204 420 206
rect 422 204 431 206
rect 417 188 431 204
rect 433 199 441 206
rect 433 197 436 199
rect 438 197 441 199
rect 433 192 441 197
rect 433 190 436 192
rect 438 190 441 192
rect 433 188 441 190
rect 443 199 451 206
rect 443 197 446 199
rect 448 197 451 199
rect 443 188 451 197
rect 453 209 458 215
rect 474 213 481 215
rect 474 211 476 213
rect 478 211 481 213
rect 453 207 460 209
rect 453 205 456 207
rect 458 205 460 207
rect 453 203 460 205
rect 453 188 458 203
rect 474 203 481 211
rect 475 199 481 203
rect 483 199 488 215
rect 490 203 498 215
rect 490 201 493 203
rect 495 201 498 203
rect 490 199 498 201
rect 500 199 505 215
rect 507 213 515 215
rect 507 211 510 213
rect 512 211 515 213
rect 507 199 515 211
rect 475 195 479 199
rect 466 193 471 195
rect 464 191 471 193
rect 464 189 466 191
rect 468 189 471 191
rect 464 187 471 189
rect 473 187 479 195
rect 510 197 515 199
rect 517 208 522 215
rect 538 213 545 215
rect 538 211 540 213
rect 542 211 545 213
rect 517 206 524 208
rect 517 204 520 206
rect 522 204 524 206
rect 517 202 524 204
rect 538 203 545 211
rect 517 197 522 202
rect 539 199 545 203
rect 547 199 552 215
rect 554 203 562 215
rect 554 201 557 203
rect 559 201 562 203
rect 554 199 562 201
rect 564 199 569 215
rect 571 213 579 215
rect 571 211 574 213
rect 576 211 579 213
rect 571 199 579 211
rect 539 195 543 199
rect 530 193 535 195
rect 528 191 535 193
rect 528 189 530 191
rect 532 189 535 191
rect 528 187 535 189
rect 537 187 543 195
rect 574 197 579 199
rect 581 208 586 215
rect 602 213 609 215
rect 602 211 604 213
rect 606 211 609 213
rect 581 206 588 208
rect 581 204 584 206
rect 586 204 588 206
rect 581 202 588 204
rect 602 203 609 211
rect 581 197 586 202
rect 603 199 609 203
rect 611 199 616 215
rect 618 203 626 215
rect 618 201 621 203
rect 623 201 626 203
rect 618 199 626 201
rect 628 199 633 215
rect 635 213 643 215
rect 635 211 638 213
rect 640 211 643 213
rect 635 199 643 211
rect 603 195 607 199
rect 594 193 599 195
rect 592 191 599 193
rect 592 189 594 191
rect 596 189 599 191
rect 592 187 599 189
rect 601 187 607 195
rect 638 197 643 199
rect 645 208 650 215
rect 645 206 652 208
rect 645 204 648 206
rect 650 204 652 206
rect 645 202 652 204
rect 645 197 650 202
rect 9 95 14 110
rect 7 93 14 95
rect 7 91 9 93
rect 11 91 14 93
rect 7 89 14 91
rect 9 83 14 89
rect 16 101 24 110
rect 16 99 19 101
rect 21 99 24 101
rect 16 92 24 99
rect 26 108 34 110
rect 26 106 29 108
rect 31 106 34 108
rect 26 101 34 106
rect 26 99 29 101
rect 31 99 34 101
rect 26 92 34 99
rect 36 94 50 110
rect 36 92 45 94
rect 47 92 50 94
rect 16 83 21 92
rect 38 87 50 92
rect 38 85 45 87
rect 47 85 50 87
rect 38 83 50 85
rect 52 108 59 110
rect 52 106 55 108
rect 57 106 59 108
rect 52 104 59 106
rect 52 83 57 104
rect 92 103 98 110
rect 71 94 78 103
rect 71 92 73 94
rect 75 92 78 94
rect 71 90 78 92
rect 80 101 88 103
rect 80 99 83 101
rect 85 99 88 101
rect 80 94 88 99
rect 80 92 83 94
rect 85 92 88 94
rect 80 90 88 92
rect 90 96 98 103
rect 90 94 93 96
rect 95 94 98 96
rect 90 92 98 94
rect 100 108 107 110
rect 100 106 103 108
rect 105 106 107 108
rect 100 101 107 106
rect 100 99 103 101
rect 105 99 107 101
rect 100 97 107 99
rect 100 92 105 97
rect 113 95 118 110
rect 111 93 118 95
rect 90 90 96 92
rect 111 91 113 93
rect 115 91 118 93
rect 111 89 118 91
rect 113 83 118 89
rect 120 101 128 110
rect 120 99 123 101
rect 125 99 128 101
rect 120 92 128 99
rect 130 108 138 110
rect 130 106 133 108
rect 135 106 138 108
rect 130 101 138 106
rect 130 99 133 101
rect 135 99 138 101
rect 130 92 138 99
rect 140 94 154 110
rect 140 92 149 94
rect 151 92 154 94
rect 120 83 125 92
rect 142 87 154 92
rect 142 85 149 87
rect 151 85 154 87
rect 142 83 154 85
rect 156 108 163 110
rect 156 106 159 108
rect 161 106 163 108
rect 156 104 163 106
rect 156 83 161 104
rect 196 103 202 110
rect 175 94 182 103
rect 175 92 177 94
rect 179 92 182 94
rect 175 90 182 92
rect 184 101 192 103
rect 184 99 187 101
rect 189 99 192 101
rect 184 94 192 99
rect 184 92 187 94
rect 189 92 192 94
rect 184 90 192 92
rect 194 96 202 103
rect 194 94 197 96
rect 199 94 202 96
rect 194 92 202 94
rect 204 108 211 110
rect 204 106 207 108
rect 209 106 211 108
rect 204 101 211 106
rect 234 104 242 111
rect 204 99 207 101
rect 209 99 211 101
rect 204 97 211 99
rect 204 92 209 97
rect 217 96 222 104
rect 215 94 222 96
rect 215 92 217 94
rect 219 92 222 94
rect 194 90 200 92
rect 215 90 222 92
rect 217 83 222 90
rect 224 83 229 104
rect 231 93 242 104
rect 244 106 249 111
rect 244 104 251 106
rect 244 102 247 104
rect 249 102 251 104
rect 244 97 251 102
rect 244 95 247 97
rect 249 95 251 97
rect 258 95 263 110
rect 244 93 251 95
rect 256 93 263 95
rect 231 87 240 93
rect 256 91 258 93
rect 260 91 263 93
rect 256 89 263 91
rect 231 85 236 87
rect 238 85 240 87
rect 231 83 240 85
rect 258 83 263 89
rect 265 101 273 110
rect 265 99 268 101
rect 270 99 273 101
rect 265 92 273 99
rect 275 108 283 110
rect 275 106 278 108
rect 280 106 283 108
rect 275 101 283 106
rect 275 99 278 101
rect 280 99 283 101
rect 275 92 283 99
rect 285 94 299 110
rect 285 92 294 94
rect 296 92 299 94
rect 265 83 270 92
rect 287 87 299 92
rect 287 85 294 87
rect 296 85 299 87
rect 287 83 299 85
rect 301 108 308 110
rect 301 106 304 108
rect 306 106 308 108
rect 301 104 308 106
rect 301 83 306 104
rect 341 103 347 110
rect 320 94 327 103
rect 320 92 322 94
rect 324 92 327 94
rect 320 90 327 92
rect 329 101 337 103
rect 329 99 332 101
rect 334 99 337 101
rect 329 94 337 99
rect 329 92 332 94
rect 334 92 337 94
rect 329 90 337 92
rect 339 96 347 103
rect 339 94 342 96
rect 344 94 347 96
rect 339 92 347 94
rect 349 108 356 110
rect 349 106 352 108
rect 354 106 356 108
rect 349 101 356 106
rect 379 104 387 111
rect 349 99 352 101
rect 354 99 356 101
rect 349 97 356 99
rect 349 92 354 97
rect 362 96 367 104
rect 360 94 367 96
rect 360 92 362 94
rect 364 92 367 94
rect 339 90 345 92
rect 360 90 367 92
rect 362 83 367 90
rect 369 83 374 104
rect 376 93 387 104
rect 389 106 394 111
rect 408 108 415 110
rect 408 106 410 108
rect 412 106 415 108
rect 389 104 396 106
rect 408 104 415 106
rect 389 102 392 104
rect 394 102 396 104
rect 389 97 396 102
rect 389 95 392 97
rect 394 95 396 97
rect 389 93 396 95
rect 376 87 385 93
rect 376 85 381 87
rect 383 85 385 87
rect 376 83 385 85
rect 410 83 415 104
rect 417 94 431 110
rect 417 92 420 94
rect 422 92 431 94
rect 433 108 441 110
rect 433 106 436 108
rect 438 106 441 108
rect 433 101 441 106
rect 433 99 436 101
rect 438 99 441 101
rect 433 92 441 99
rect 443 101 451 110
rect 443 99 446 101
rect 448 99 451 101
rect 443 92 451 99
rect 417 87 429 92
rect 417 85 420 87
rect 422 85 429 87
rect 417 83 429 85
rect 446 83 451 92
rect 453 95 458 110
rect 464 109 471 111
rect 464 107 466 109
rect 468 107 471 109
rect 464 105 471 107
rect 466 103 471 105
rect 473 103 479 111
rect 475 99 479 103
rect 528 109 535 111
rect 528 107 530 109
rect 532 107 535 109
rect 528 105 535 107
rect 530 103 535 105
rect 537 103 543 111
rect 510 99 515 101
rect 453 93 460 95
rect 475 95 481 99
rect 453 91 456 93
rect 458 91 460 93
rect 453 89 460 91
rect 453 83 458 89
rect 474 87 481 95
rect 474 85 476 87
rect 478 85 481 87
rect 474 83 481 85
rect 483 83 488 99
rect 490 97 498 99
rect 490 95 493 97
rect 495 95 498 97
rect 490 83 498 95
rect 500 83 505 99
rect 507 87 515 99
rect 507 85 510 87
rect 512 85 515 87
rect 507 83 515 85
rect 517 96 522 101
rect 539 99 543 103
rect 592 109 599 111
rect 592 107 594 109
rect 596 107 599 109
rect 592 105 599 107
rect 594 103 599 105
rect 601 103 607 111
rect 574 99 579 101
rect 517 94 524 96
rect 539 95 545 99
rect 517 92 520 94
rect 522 92 524 94
rect 517 90 524 92
rect 517 83 522 90
rect 538 87 545 95
rect 538 85 540 87
rect 542 85 545 87
rect 538 83 545 85
rect 547 83 552 99
rect 554 97 562 99
rect 554 95 557 97
rect 559 95 562 97
rect 554 83 562 95
rect 564 83 569 99
rect 571 87 579 99
rect 571 85 574 87
rect 576 85 579 87
rect 571 83 579 85
rect 581 96 586 101
rect 603 99 607 103
rect 638 99 643 101
rect 581 94 588 96
rect 603 95 609 99
rect 581 92 584 94
rect 586 92 588 94
rect 581 90 588 92
rect 581 83 586 90
rect 602 87 609 95
rect 602 85 604 87
rect 606 85 609 87
rect 602 83 609 85
rect 611 83 616 99
rect 618 97 626 99
rect 618 95 621 97
rect 623 95 626 97
rect 618 83 626 95
rect 628 83 633 99
rect 635 87 643 99
rect 635 85 638 87
rect 640 85 643 87
rect 635 83 643 85
rect 645 96 650 101
rect 645 94 652 96
rect 645 92 648 94
rect 650 92 652 94
rect 645 90 652 92
rect 645 83 650 90
rect 18 69 27 71
rect 18 67 20 69
rect 22 67 27 69
rect 18 61 27 67
rect 7 59 14 61
rect 7 57 9 59
rect 11 57 14 59
rect 7 52 14 57
rect 7 50 9 52
rect 11 50 14 52
rect 7 48 14 50
rect 9 43 14 48
rect 16 50 27 61
rect 29 50 34 71
rect 36 64 41 71
rect 36 62 43 64
rect 58 62 64 64
rect 36 60 39 62
rect 41 60 43 62
rect 36 58 43 60
rect 36 50 41 58
rect 49 57 54 62
rect 47 55 54 57
rect 47 53 49 55
rect 51 53 54 55
rect 16 43 24 50
rect 47 48 54 53
rect 47 46 49 48
rect 51 46 54 48
rect 47 44 54 46
rect 56 60 64 62
rect 56 58 59 60
rect 61 58 64 60
rect 56 51 64 58
rect 66 62 74 64
rect 66 60 69 62
rect 71 60 74 62
rect 66 55 74 60
rect 66 53 69 55
rect 71 53 74 55
rect 66 51 74 53
rect 76 62 83 64
rect 76 60 79 62
rect 81 60 83 62
rect 76 51 83 60
rect 56 44 62 51
rect 97 50 102 71
rect 95 48 102 50
rect 95 46 97 48
rect 99 46 102 48
rect 95 44 102 46
rect 104 69 116 71
rect 104 67 107 69
rect 109 67 116 69
rect 104 62 116 67
rect 133 62 138 71
rect 104 60 107 62
rect 109 60 118 62
rect 104 44 118 60
rect 120 55 128 62
rect 120 53 123 55
rect 125 53 128 55
rect 120 48 128 53
rect 120 46 123 48
rect 125 46 128 48
rect 120 44 128 46
rect 130 55 138 62
rect 130 53 133 55
rect 135 53 138 55
rect 130 44 138 53
rect 140 65 145 71
rect 140 63 147 65
rect 140 61 143 63
rect 145 61 147 63
rect 162 62 168 64
rect 140 59 147 61
rect 140 44 145 59
rect 153 57 158 62
rect 151 55 158 57
rect 151 53 153 55
rect 155 53 158 55
rect 151 48 158 53
rect 151 46 153 48
rect 155 46 158 48
rect 151 44 158 46
rect 160 60 168 62
rect 160 58 163 60
rect 165 58 168 60
rect 160 51 168 58
rect 170 62 178 64
rect 170 60 173 62
rect 175 60 178 62
rect 170 55 178 60
rect 170 53 173 55
rect 175 53 178 55
rect 170 51 178 53
rect 180 62 187 64
rect 180 60 183 62
rect 185 60 187 62
rect 180 51 187 60
rect 160 44 166 51
rect 201 50 206 71
rect 199 48 206 50
rect 199 46 201 48
rect 203 46 206 48
rect 199 44 206 46
rect 208 69 220 71
rect 208 67 211 69
rect 213 67 220 69
rect 208 62 220 67
rect 237 62 242 71
rect 208 60 211 62
rect 213 60 222 62
rect 208 44 222 60
rect 224 55 232 62
rect 224 53 227 55
rect 229 53 232 55
rect 224 48 232 53
rect 224 46 227 48
rect 229 46 232 48
rect 224 44 232 46
rect 234 55 242 62
rect 234 53 237 55
rect 239 53 242 55
rect 234 44 242 53
rect 244 65 249 71
rect 258 65 263 71
rect 244 63 251 65
rect 244 61 247 63
rect 249 61 251 63
rect 244 59 251 61
rect 256 63 263 65
rect 256 61 258 63
rect 260 61 263 63
rect 256 59 263 61
rect 244 44 249 59
rect 258 44 263 59
rect 265 62 270 71
rect 287 69 299 71
rect 287 67 294 69
rect 296 67 299 69
rect 287 62 299 67
rect 265 55 273 62
rect 265 53 268 55
rect 270 53 273 55
rect 265 44 273 53
rect 275 55 283 62
rect 275 53 278 55
rect 280 53 283 55
rect 275 48 283 53
rect 275 46 278 48
rect 280 46 283 48
rect 275 44 283 46
rect 285 60 294 62
rect 296 60 299 62
rect 285 44 299 60
rect 301 50 306 71
rect 320 62 327 64
rect 320 60 322 62
rect 324 60 327 62
rect 320 51 327 60
rect 329 62 337 64
rect 329 60 332 62
rect 334 60 337 62
rect 329 55 337 60
rect 329 53 332 55
rect 334 53 337 55
rect 329 51 337 53
rect 339 62 345 64
rect 362 64 367 71
rect 360 62 367 64
rect 339 60 347 62
rect 339 58 342 60
rect 344 58 347 60
rect 339 51 347 58
rect 301 48 308 50
rect 301 46 304 48
rect 306 46 308 48
rect 301 44 308 46
rect 341 44 347 51
rect 349 57 354 62
rect 360 60 362 62
rect 364 60 367 62
rect 360 58 367 60
rect 349 55 356 57
rect 349 53 352 55
rect 354 53 356 55
rect 349 48 356 53
rect 362 50 367 58
rect 369 50 374 71
rect 376 69 385 71
rect 376 67 381 69
rect 383 67 385 69
rect 376 61 385 67
rect 376 50 387 61
rect 349 46 352 48
rect 354 46 356 48
rect 349 44 356 46
rect 379 43 387 50
rect 389 59 396 61
rect 389 57 392 59
rect 394 57 396 59
rect 389 52 396 57
rect 389 50 392 52
rect 394 50 396 52
rect 410 50 415 71
rect 389 48 396 50
rect 408 48 415 50
rect 389 43 394 48
rect 408 46 410 48
rect 412 46 415 48
rect 408 44 415 46
rect 417 69 429 71
rect 417 67 420 69
rect 422 67 429 69
rect 417 62 429 67
rect 446 62 451 71
rect 417 60 420 62
rect 422 60 431 62
rect 417 44 431 60
rect 433 55 441 62
rect 433 53 436 55
rect 438 53 441 55
rect 433 48 441 53
rect 433 46 436 48
rect 438 46 441 48
rect 433 44 441 46
rect 443 55 451 62
rect 443 53 446 55
rect 448 53 451 55
rect 443 44 451 53
rect 453 65 458 71
rect 474 69 481 71
rect 474 67 476 69
rect 478 67 481 69
rect 453 63 460 65
rect 453 61 456 63
rect 458 61 460 63
rect 453 59 460 61
rect 453 44 458 59
rect 474 59 481 67
rect 475 55 481 59
rect 483 55 488 71
rect 490 59 498 71
rect 490 57 493 59
rect 495 57 498 59
rect 490 55 498 57
rect 500 55 505 71
rect 507 69 515 71
rect 507 67 510 69
rect 512 67 515 69
rect 507 55 515 67
rect 475 51 479 55
rect 466 49 471 51
rect 464 47 471 49
rect 464 45 466 47
rect 468 45 471 47
rect 464 43 471 45
rect 473 43 479 51
rect 510 53 515 55
rect 517 64 522 71
rect 538 69 545 71
rect 538 67 540 69
rect 542 67 545 69
rect 517 62 524 64
rect 517 60 520 62
rect 522 60 524 62
rect 517 58 524 60
rect 538 59 545 67
rect 517 53 522 58
rect 539 55 545 59
rect 547 55 552 71
rect 554 59 562 71
rect 554 57 557 59
rect 559 57 562 59
rect 554 55 562 57
rect 564 55 569 71
rect 571 69 579 71
rect 571 67 574 69
rect 576 67 579 69
rect 571 55 579 67
rect 539 51 543 55
rect 530 49 535 51
rect 528 47 535 49
rect 528 45 530 47
rect 532 45 535 47
rect 528 43 535 45
rect 537 43 543 51
rect 574 53 579 55
rect 581 64 586 71
rect 602 69 609 71
rect 602 67 604 69
rect 606 67 609 69
rect 581 62 588 64
rect 581 60 584 62
rect 586 60 588 62
rect 581 58 588 60
rect 602 59 609 67
rect 581 53 586 58
rect 603 55 609 59
rect 611 55 616 71
rect 618 59 626 71
rect 618 57 621 59
rect 623 57 626 59
rect 618 55 626 57
rect 628 55 633 71
rect 635 69 643 71
rect 635 67 638 69
rect 640 67 643 69
rect 635 55 643 67
rect 603 51 607 55
rect 594 49 599 51
rect 592 47 599 49
rect 592 45 594 47
rect 596 45 599 47
rect 592 43 599 45
rect 601 43 607 51
rect 638 53 643 55
rect 645 64 650 71
rect 645 62 652 64
rect 645 60 648 62
rect 650 60 652 62
rect 645 58 652 60
rect 645 53 650 58
<< alu1 >>
rect 3 578 656 581
rect 3 576 4 578
rect 6 576 656 578
rect 3 574 9 576
rect 11 574 62 576
rect 64 574 92 576
rect 94 574 102 576
rect 104 574 113 576
rect 115 574 166 576
rect 168 574 196 576
rect 198 574 206 576
rect 208 574 246 576
rect 248 574 258 576
rect 260 574 311 576
rect 313 574 341 576
rect 343 574 351 576
rect 353 574 391 576
rect 393 574 403 576
rect 405 574 456 576
rect 458 574 656 576
rect 3 573 656 574
rect 7 566 31 567
rect 7 564 27 566
rect 29 564 31 566
rect 7 563 31 564
rect 7 535 11 563
rect 46 559 59 560
rect 46 557 55 559
rect 57 557 59 559
rect 46 555 59 557
rect 46 553 47 555
rect 49 554 59 555
rect 49 553 51 554
rect 7 533 23 535
rect 7 531 19 533
rect 21 531 23 533
rect 7 530 23 531
rect 46 546 51 553
rect 78 559 83 560
rect 78 557 80 559
rect 82 557 83 559
rect 78 551 83 557
rect 95 564 107 568
rect 95 562 103 564
rect 105 562 107 564
rect 78 550 92 551
rect 78 548 86 550
rect 88 548 89 550
rect 91 548 92 550
rect 78 547 92 548
rect 62 542 67 544
rect 62 540 63 542
rect 65 540 67 542
rect 62 535 67 540
rect 62 533 63 535
rect 65 533 67 535
rect 62 528 67 533
rect 71 542 84 543
rect 71 540 76 542
rect 78 540 81 542
rect 83 540 84 542
rect 71 539 84 540
rect 71 535 75 539
rect 103 550 107 562
rect 103 548 104 550
rect 106 548 107 550
rect 103 542 107 548
rect 71 533 72 535
rect 74 533 75 535
rect 71 530 75 533
rect 102 540 107 542
rect 102 538 103 540
rect 105 538 107 540
rect 102 533 107 538
rect 55 522 67 528
rect 102 531 103 533
rect 105 531 107 533
rect 102 529 107 531
rect 111 566 135 567
rect 111 564 131 566
rect 133 564 135 566
rect 111 563 135 564
rect 111 542 115 563
rect 150 559 163 560
rect 150 557 159 559
rect 161 557 163 559
rect 150 555 163 557
rect 150 553 151 555
rect 153 554 163 555
rect 153 553 155 554
rect 111 540 112 542
rect 114 540 115 542
rect 111 535 115 540
rect 111 533 127 535
rect 111 531 123 533
rect 125 531 127 533
rect 111 530 127 531
rect 150 546 155 553
rect 182 559 187 560
rect 182 557 184 559
rect 186 557 187 559
rect 182 551 187 557
rect 199 564 211 568
rect 344 567 356 568
rect 199 562 207 564
rect 209 562 211 564
rect 182 550 196 551
rect 182 548 190 550
rect 192 548 196 550
rect 182 547 196 548
rect 166 542 171 544
rect 166 540 167 542
rect 169 540 171 542
rect 166 535 171 540
rect 166 533 167 535
rect 169 533 171 535
rect 166 528 171 533
rect 175 542 188 543
rect 175 540 180 542
rect 182 540 188 542
rect 175 539 188 540
rect 175 535 179 539
rect 207 542 211 562
rect 256 566 280 567
rect 256 564 276 566
rect 278 564 280 566
rect 256 563 280 564
rect 215 551 219 560
rect 215 550 236 551
rect 215 548 216 550
rect 218 548 230 550
rect 232 548 236 550
rect 215 547 236 548
rect 246 559 251 561
rect 246 557 247 559
rect 249 557 251 559
rect 246 555 251 557
rect 175 533 176 535
rect 178 533 179 535
rect 175 530 179 533
rect 206 540 211 542
rect 206 538 207 540
rect 209 538 211 540
rect 206 537 211 538
rect 206 535 208 537
rect 210 535 211 537
rect 206 533 211 535
rect 159 522 171 528
rect 206 531 207 533
rect 209 531 211 533
rect 206 529 211 531
rect 215 541 220 543
rect 222 541 236 543
rect 215 539 236 541
rect 215 537 219 539
rect 215 535 216 537
rect 218 535 219 537
rect 215 530 219 535
rect 247 536 251 555
rect 249 534 251 536
rect 247 529 251 534
rect 256 535 260 563
rect 295 558 308 560
rect 295 556 303 558
rect 305 556 308 558
rect 295 555 308 556
rect 295 553 296 555
rect 298 554 308 555
rect 298 553 300 554
rect 256 533 272 535
rect 256 531 257 533
rect 259 531 268 533
rect 270 531 272 533
rect 256 530 272 531
rect 295 546 300 553
rect 327 558 332 560
rect 327 556 329 558
rect 331 556 332 558
rect 327 551 332 556
rect 344 565 353 567
rect 355 565 356 567
rect 344 564 356 565
rect 436 566 460 567
rect 344 562 352 564
rect 354 562 356 564
rect 327 550 341 551
rect 327 548 335 550
rect 337 548 341 550
rect 327 547 341 548
rect 311 542 316 544
rect 311 540 312 542
rect 314 540 316 542
rect 249 527 251 529
rect 238 523 251 527
rect 311 534 316 540
rect 311 532 313 534
rect 315 532 316 534
rect 311 528 316 532
rect 320 542 333 543
rect 320 540 325 542
rect 327 540 333 542
rect 320 539 333 540
rect 320 534 324 539
rect 352 542 356 562
rect 436 564 438 566
rect 440 564 460 566
rect 436 563 460 564
rect 360 558 364 560
rect 360 556 361 558
rect 363 556 364 558
rect 360 551 364 556
rect 360 550 381 551
rect 360 548 375 550
rect 377 548 381 550
rect 360 547 381 548
rect 391 559 396 561
rect 391 557 392 559
rect 394 557 396 559
rect 391 555 396 557
rect 320 532 321 534
rect 323 532 324 534
rect 320 530 324 532
rect 351 540 356 542
rect 351 538 352 540
rect 354 538 356 540
rect 351 533 356 538
rect 247 522 251 523
rect 304 522 316 528
rect 351 531 352 533
rect 354 531 356 533
rect 351 529 356 531
rect 360 541 365 543
rect 367 541 381 543
rect 360 539 381 541
rect 360 533 364 539
rect 392 543 396 555
rect 408 558 421 560
rect 408 556 411 558
rect 413 556 421 558
rect 408 555 421 556
rect 408 554 418 555
rect 416 553 418 554
rect 420 553 421 555
rect 392 541 393 543
rect 395 541 396 543
rect 360 531 361 533
rect 363 531 364 533
rect 360 530 364 531
rect 392 536 396 541
rect 394 534 396 536
rect 392 529 396 534
rect 394 527 396 529
rect 383 523 396 527
rect 392 522 396 523
rect 400 542 405 544
rect 400 540 402 542
rect 404 540 405 542
rect 400 533 405 540
rect 416 546 421 553
rect 456 558 460 563
rect 456 556 457 558
rect 459 556 460 558
rect 400 531 402 533
rect 404 531 405 533
rect 400 528 405 531
rect 400 522 412 528
rect 456 535 460 556
rect 520 566 524 568
rect 519 564 524 566
rect 519 562 520 564
rect 522 562 524 564
rect 519 560 524 562
rect 471 558 484 559
rect 471 556 472 558
rect 474 556 484 558
rect 471 555 484 556
rect 478 550 484 555
rect 478 548 479 550
rect 481 548 484 550
rect 478 546 484 548
rect 504 545 508 552
rect 504 544 506 545
rect 496 543 506 544
rect 496 541 497 543
rect 499 541 508 543
rect 496 538 508 541
rect 444 533 460 535
rect 444 531 446 533
rect 448 531 460 533
rect 444 530 460 531
rect 464 531 477 535
rect 464 530 469 531
rect 520 534 524 560
rect 584 566 588 568
rect 583 564 588 566
rect 583 562 584 564
rect 586 562 588 564
rect 583 560 588 562
rect 535 558 548 559
rect 535 556 536 558
rect 538 556 548 558
rect 535 555 548 556
rect 542 550 548 555
rect 542 548 543 550
rect 545 548 548 550
rect 542 546 548 548
rect 584 558 588 560
rect 568 545 572 552
rect 584 556 585 558
rect 587 556 588 558
rect 568 544 570 545
rect 560 543 570 544
rect 560 541 561 543
rect 563 541 572 543
rect 560 538 572 541
rect 520 532 521 534
rect 523 532 524 534
rect 464 528 466 530
rect 468 528 469 530
rect 464 525 469 528
rect 520 527 524 532
rect 511 526 524 527
rect 464 523 466 525
rect 468 523 469 525
rect 511 524 520 526
rect 522 524 524 526
rect 511 523 524 524
rect 528 531 541 535
rect 528 530 533 531
rect 528 528 530 530
rect 532 528 533 530
rect 528 525 533 528
rect 584 527 588 556
rect 648 566 652 568
rect 647 564 652 566
rect 647 562 648 564
rect 650 562 652 564
rect 647 560 652 562
rect 599 558 612 559
rect 599 556 600 558
rect 602 556 612 558
rect 599 555 612 556
rect 606 550 612 555
rect 606 548 607 550
rect 609 548 612 550
rect 606 546 612 548
rect 632 545 636 552
rect 632 544 634 545
rect 624 543 634 544
rect 624 541 636 543
rect 624 539 625 541
rect 627 539 636 541
rect 624 538 636 539
rect 575 526 588 527
rect 528 523 530 525
rect 532 523 533 525
rect 575 524 584 526
rect 586 524 588 526
rect 575 523 588 524
rect 592 531 605 535
rect 592 530 597 531
rect 592 528 594 530
rect 596 528 597 530
rect 592 525 597 528
rect 648 527 652 560
rect 639 526 652 527
rect 592 523 594 525
rect 596 523 597 525
rect 639 524 648 526
rect 650 524 652 526
rect 639 523 652 524
rect 464 522 469 523
rect 528 522 533 523
rect 592 522 597 523
rect 3 516 656 517
rect 3 514 29 516
rect 31 514 102 516
rect 104 514 133 516
rect 135 514 206 516
rect 208 514 246 516
rect 248 514 278 516
rect 280 514 351 516
rect 353 514 391 516
rect 393 514 436 516
rect 438 514 656 516
rect 3 505 656 514
rect 3 504 252 505
rect 3 502 10 504
rect 12 502 50 504
rect 52 502 123 504
rect 125 502 154 504
rect 156 502 227 504
rect 229 503 252 504
rect 254 504 656 505
rect 254 503 278 504
rect 229 502 278 503
rect 280 502 351 504
rect 353 502 391 504
rect 393 502 436 504
rect 438 502 656 504
rect 3 501 656 502
rect 7 495 11 496
rect 7 491 20 495
rect 7 489 9 491
rect 7 484 11 489
rect 7 482 9 484
rect 7 472 11 482
rect 39 483 43 488
rect 7 470 8 472
rect 10 470 11 472
rect 7 463 11 470
rect 39 481 40 483
rect 42 481 43 483
rect 39 479 43 481
rect 22 477 43 479
rect 22 475 36 477
rect 38 475 43 477
rect 47 487 52 489
rect 47 485 49 487
rect 51 485 52 487
rect 87 490 99 496
rect 47 483 52 485
rect 47 481 48 483
rect 50 481 52 483
rect 47 480 52 481
rect 47 478 49 480
rect 51 478 52 480
rect 47 476 52 478
rect 79 485 83 488
rect 79 483 80 485
rect 82 483 83 485
rect 7 461 12 463
rect 7 459 9 461
rect 11 459 12 461
rect 7 457 12 459
rect 22 470 43 471
rect 22 468 26 470
rect 28 468 40 470
rect 42 468 43 470
rect 22 467 43 468
rect 39 458 43 467
rect 47 456 51 476
rect 79 479 83 483
rect 70 478 83 479
rect 70 476 76 478
rect 78 476 83 478
rect 70 475 83 476
rect 87 485 92 490
rect 87 483 89 485
rect 91 483 92 485
rect 87 478 92 483
rect 87 476 89 478
rect 91 476 92 478
rect 87 474 92 476
rect 62 470 76 471
rect 62 468 66 470
rect 68 468 76 470
rect 62 467 76 468
rect 47 454 49 456
rect 51 454 59 456
rect 47 450 59 454
rect 71 461 76 467
rect 71 459 72 461
rect 74 459 76 461
rect 71 458 76 459
rect 103 465 108 472
rect 131 487 147 488
rect 131 485 133 487
rect 135 485 147 487
rect 131 483 147 485
rect 143 478 147 483
rect 143 476 144 478
rect 146 476 147 478
rect 103 464 105 465
rect 95 463 105 464
rect 107 463 108 465
rect 95 461 108 463
rect 95 459 97 461
rect 99 459 108 461
rect 95 458 108 459
rect 143 455 147 476
rect 123 454 147 455
rect 123 452 125 454
rect 127 452 147 454
rect 123 451 147 452
rect 151 487 156 489
rect 151 485 153 487
rect 155 485 156 487
rect 191 490 203 496
rect 151 480 156 485
rect 151 478 153 480
rect 155 478 156 480
rect 151 476 156 478
rect 183 485 187 488
rect 183 483 184 485
rect 186 483 187 485
rect 151 470 155 476
rect 151 468 152 470
rect 154 468 155 470
rect 151 456 155 468
rect 183 479 187 483
rect 174 478 187 479
rect 174 476 175 478
rect 177 476 180 478
rect 182 476 187 478
rect 174 475 187 476
rect 191 485 196 490
rect 191 483 193 485
rect 195 483 196 485
rect 191 478 196 483
rect 191 476 193 478
rect 195 476 196 478
rect 191 474 196 476
rect 166 470 180 471
rect 166 468 170 470
rect 172 468 177 470
rect 179 468 180 470
rect 166 467 180 468
rect 151 454 153 456
rect 155 454 163 456
rect 151 450 163 454
rect 175 461 180 467
rect 175 459 176 461
rect 178 459 180 461
rect 175 458 180 459
rect 207 465 212 472
rect 235 487 251 488
rect 235 485 237 487
rect 239 486 251 487
rect 239 485 243 486
rect 235 484 243 485
rect 245 484 251 486
rect 235 483 251 484
rect 207 464 209 465
rect 199 463 209 464
rect 211 463 212 465
rect 199 461 212 463
rect 199 459 201 461
rect 203 459 212 461
rect 199 458 212 459
rect 247 455 251 483
rect 227 454 251 455
rect 227 452 229 454
rect 231 452 251 454
rect 227 451 251 452
rect 256 487 272 488
rect 256 486 268 487
rect 256 484 257 486
rect 259 485 268 486
rect 270 485 272 487
rect 259 484 272 485
rect 256 483 272 484
rect 256 455 260 483
rect 304 490 316 496
rect 311 487 316 490
rect 311 485 313 487
rect 315 485 316 487
rect 295 465 300 472
rect 311 478 316 485
rect 311 476 312 478
rect 314 476 316 478
rect 311 474 316 476
rect 320 487 324 488
rect 320 485 321 487
rect 323 485 324 487
rect 320 479 324 485
rect 392 495 396 496
rect 383 491 396 495
rect 351 487 356 489
rect 320 478 333 479
rect 320 476 325 478
rect 327 476 333 478
rect 320 475 333 476
rect 295 463 296 465
rect 298 464 300 465
rect 298 463 308 464
rect 295 462 308 463
rect 295 460 303 462
rect 305 460 308 462
rect 295 458 308 460
rect 327 470 341 471
rect 327 468 335 470
rect 337 468 341 470
rect 327 467 341 468
rect 351 485 352 487
rect 354 485 356 487
rect 351 480 356 485
rect 351 478 352 480
rect 354 478 356 480
rect 351 476 356 478
rect 327 461 332 467
rect 327 459 329 461
rect 331 459 332 461
rect 327 458 332 459
rect 256 454 280 455
rect 256 452 276 454
rect 278 452 280 454
rect 352 456 356 476
rect 360 487 364 488
rect 360 485 361 487
rect 363 485 364 487
rect 360 479 364 485
rect 360 477 381 479
rect 360 475 365 477
rect 367 475 381 477
rect 360 470 381 471
rect 360 468 375 470
rect 377 468 381 470
rect 360 467 381 468
rect 394 489 396 491
rect 392 484 396 489
rect 394 482 396 484
rect 360 461 364 467
rect 392 477 396 482
rect 392 475 393 477
rect 395 475 396 477
rect 392 463 396 475
rect 400 490 412 496
rect 464 495 469 496
rect 528 495 533 496
rect 592 495 597 496
rect 464 493 465 495
rect 467 493 469 495
rect 400 487 405 490
rect 400 485 402 487
rect 404 485 405 487
rect 400 478 405 485
rect 464 490 469 493
rect 511 494 524 495
rect 511 492 520 494
rect 522 492 524 494
rect 400 476 402 478
rect 404 476 405 478
rect 400 474 405 476
rect 360 459 361 461
rect 363 459 364 461
rect 360 458 364 459
rect 391 461 396 463
rect 391 459 392 461
rect 394 459 396 461
rect 391 457 396 459
rect 416 465 421 472
rect 464 488 466 490
rect 468 488 469 490
rect 511 491 524 492
rect 444 487 460 488
rect 444 485 446 487
rect 448 485 460 487
rect 444 483 460 485
rect 464 487 469 488
rect 464 483 477 487
rect 416 464 418 465
rect 408 463 418 464
rect 420 463 421 465
rect 408 461 421 463
rect 408 459 411 461
rect 413 459 421 461
rect 408 458 421 459
rect 456 462 460 483
rect 456 460 457 462
rect 459 460 460 462
rect 256 451 280 452
rect 344 454 352 456
rect 354 454 356 456
rect 456 455 460 460
rect 344 453 356 454
rect 344 451 353 453
rect 355 451 356 453
rect 344 450 356 451
rect 436 454 460 455
rect 436 452 438 454
rect 440 452 460 454
rect 478 470 484 472
rect 478 468 479 470
rect 481 468 484 470
rect 478 463 484 468
rect 471 462 484 463
rect 471 460 472 462
rect 474 460 484 462
rect 496 477 508 480
rect 496 475 497 477
rect 499 475 508 477
rect 496 474 506 475
rect 504 473 506 474
rect 504 466 508 473
rect 520 486 524 491
rect 520 484 521 486
rect 523 484 524 486
rect 471 459 484 460
rect 520 458 524 484
rect 528 493 530 495
rect 532 493 533 495
rect 528 490 533 493
rect 575 494 588 495
rect 575 492 584 494
rect 586 492 588 494
rect 528 488 530 490
rect 532 488 533 490
rect 575 491 588 492
rect 528 487 533 488
rect 528 483 541 487
rect 519 456 524 458
rect 436 451 460 452
rect 519 454 520 456
rect 522 454 524 456
rect 519 452 524 454
rect 542 470 548 472
rect 542 468 543 470
rect 545 468 548 470
rect 542 463 548 468
rect 535 462 548 463
rect 535 460 536 462
rect 538 460 548 462
rect 560 477 572 480
rect 560 475 561 477
rect 563 475 572 477
rect 560 474 570 475
rect 568 473 570 474
rect 568 466 572 473
rect 584 462 588 491
rect 592 493 594 495
rect 596 493 597 495
rect 592 490 597 493
rect 639 494 652 495
rect 639 492 648 494
rect 650 492 652 494
rect 592 488 594 490
rect 596 488 597 490
rect 639 491 652 492
rect 592 487 597 488
rect 592 483 605 487
rect 535 459 548 460
rect 584 460 585 462
rect 587 460 588 462
rect 584 458 588 460
rect 583 456 588 458
rect 520 450 524 452
rect 583 454 584 456
rect 586 454 588 456
rect 583 452 588 454
rect 606 470 612 472
rect 606 468 607 470
rect 609 468 612 470
rect 606 463 612 468
rect 599 462 612 463
rect 599 460 600 462
rect 602 460 612 462
rect 624 479 636 480
rect 624 477 625 479
rect 627 477 636 479
rect 624 475 636 477
rect 624 474 634 475
rect 632 473 634 474
rect 632 466 636 473
rect 599 459 612 460
rect 648 458 652 491
rect 647 456 652 458
rect 584 450 588 452
rect 647 454 648 456
rect 650 454 652 456
rect 647 452 652 454
rect 648 450 652 452
rect 3 444 656 445
rect 3 442 4 444
rect 6 442 10 444
rect 12 442 50 444
rect 52 442 60 444
rect 62 442 90 444
rect 92 442 143 444
rect 145 442 154 444
rect 156 442 164 444
rect 166 442 194 444
rect 196 442 247 444
rect 249 442 258 444
rect 260 442 311 444
rect 313 442 341 444
rect 343 442 351 444
rect 353 442 391 444
rect 393 442 403 444
rect 405 442 456 444
rect 458 442 656 444
rect 3 434 656 442
rect 3 432 4 434
rect 6 432 656 434
rect 3 430 9 432
rect 11 430 62 432
rect 64 430 92 432
rect 94 430 102 432
rect 104 430 113 432
rect 115 430 166 432
rect 168 430 196 432
rect 198 430 206 432
rect 208 430 246 432
rect 248 430 258 432
rect 260 430 311 432
rect 313 430 341 432
rect 343 430 351 432
rect 353 430 391 432
rect 393 430 403 432
rect 405 430 456 432
rect 458 430 656 432
rect 3 429 656 430
rect 7 422 31 423
rect 7 420 27 422
rect 29 420 31 422
rect 7 419 31 420
rect 7 391 11 419
rect 46 415 59 416
rect 46 413 55 415
rect 57 413 59 415
rect 46 411 59 413
rect 46 409 47 411
rect 49 410 59 411
rect 49 409 51 410
rect 7 389 23 391
rect 7 387 19 389
rect 21 387 23 389
rect 7 386 23 387
rect 46 402 51 409
rect 78 415 83 416
rect 78 413 80 415
rect 82 413 83 415
rect 78 407 83 413
rect 95 420 107 424
rect 95 418 103 420
rect 105 418 107 420
rect 78 406 92 407
rect 78 404 81 406
rect 83 404 86 406
rect 88 404 92 406
rect 78 403 92 404
rect 62 398 67 400
rect 62 396 63 398
rect 65 396 67 398
rect 62 391 67 396
rect 62 389 63 391
rect 65 389 67 391
rect 62 384 67 389
rect 71 398 84 399
rect 71 396 76 398
rect 78 396 81 398
rect 83 396 84 398
rect 71 395 84 396
rect 71 391 75 395
rect 103 406 107 418
rect 103 404 104 406
rect 106 404 107 406
rect 103 398 107 404
rect 71 389 72 391
rect 74 389 75 391
rect 71 386 75 389
rect 102 396 107 398
rect 102 394 103 396
rect 105 394 107 396
rect 102 389 107 394
rect 55 378 67 384
rect 102 387 103 389
rect 105 387 107 389
rect 102 385 107 387
rect 111 422 135 423
rect 111 420 131 422
rect 133 420 135 422
rect 111 419 135 420
rect 111 398 115 419
rect 150 415 163 416
rect 150 413 159 415
rect 161 413 163 415
rect 150 411 163 413
rect 150 409 151 411
rect 153 410 163 411
rect 153 409 155 410
rect 111 396 112 398
rect 114 396 115 398
rect 111 391 115 396
rect 111 389 127 391
rect 111 387 123 389
rect 125 387 127 389
rect 111 386 127 387
rect 150 402 155 409
rect 182 415 187 416
rect 182 413 184 415
rect 186 413 187 415
rect 182 407 187 413
rect 199 420 211 424
rect 344 423 356 424
rect 199 418 207 420
rect 209 418 211 420
rect 182 406 196 407
rect 182 404 190 406
rect 192 404 196 406
rect 182 403 196 404
rect 166 398 171 400
rect 166 396 167 398
rect 169 396 171 398
rect 166 391 171 396
rect 166 389 167 391
rect 169 389 171 391
rect 166 384 171 389
rect 175 398 188 399
rect 175 396 180 398
rect 182 396 188 398
rect 175 395 188 396
rect 175 391 179 395
rect 207 398 211 418
rect 256 422 280 423
rect 256 420 276 422
rect 278 420 280 422
rect 256 419 280 420
rect 215 407 219 416
rect 215 406 236 407
rect 215 404 216 406
rect 218 404 230 406
rect 232 404 236 406
rect 215 403 236 404
rect 246 415 251 417
rect 246 413 247 415
rect 249 413 251 415
rect 246 411 251 413
rect 175 389 176 391
rect 178 389 179 391
rect 175 386 179 389
rect 206 396 211 398
rect 206 394 207 396
rect 209 394 211 396
rect 206 393 211 394
rect 206 391 208 393
rect 210 391 211 393
rect 206 389 211 391
rect 159 378 171 384
rect 206 387 207 389
rect 209 387 211 389
rect 206 385 211 387
rect 215 397 220 399
rect 222 397 236 399
rect 215 395 236 397
rect 215 393 219 395
rect 215 391 216 393
rect 218 391 219 393
rect 247 409 251 411
rect 247 407 248 409
rect 250 407 251 409
rect 215 386 219 391
rect 247 392 251 407
rect 249 390 251 392
rect 247 385 251 390
rect 256 391 260 419
rect 295 414 308 416
rect 295 412 303 414
rect 305 412 308 414
rect 295 411 308 412
rect 295 409 296 411
rect 298 410 308 411
rect 298 409 300 410
rect 256 389 272 391
rect 256 387 257 389
rect 259 387 268 389
rect 270 387 272 389
rect 256 386 272 387
rect 295 402 300 409
rect 327 414 332 416
rect 327 412 329 414
rect 331 412 332 414
rect 327 407 332 412
rect 344 421 353 423
rect 355 421 356 423
rect 344 420 356 421
rect 436 422 460 423
rect 344 418 352 420
rect 354 418 356 420
rect 327 406 341 407
rect 327 404 335 406
rect 337 404 341 406
rect 327 403 341 404
rect 311 398 316 400
rect 311 396 312 398
rect 314 396 316 398
rect 249 383 251 385
rect 238 379 251 383
rect 311 389 316 396
rect 311 387 312 389
rect 314 387 316 389
rect 311 384 316 387
rect 320 398 333 399
rect 320 396 325 398
rect 327 396 333 398
rect 320 395 333 396
rect 320 389 324 395
rect 352 398 356 418
rect 436 420 438 422
rect 440 420 460 422
rect 436 419 460 420
rect 360 414 364 416
rect 360 412 361 414
rect 363 412 364 414
rect 360 407 364 412
rect 360 406 381 407
rect 360 404 375 406
rect 377 404 381 406
rect 360 403 381 404
rect 391 415 396 417
rect 391 413 392 415
rect 394 413 396 415
rect 391 411 396 413
rect 320 387 321 389
rect 323 387 324 389
rect 320 386 324 387
rect 351 396 356 398
rect 351 394 352 396
rect 354 394 356 396
rect 351 389 356 394
rect 247 378 251 379
rect 304 378 316 384
rect 351 387 352 389
rect 354 387 356 389
rect 351 385 356 387
rect 360 397 365 399
rect 367 397 381 399
rect 360 395 381 397
rect 360 389 364 395
rect 392 399 396 411
rect 408 414 421 416
rect 408 412 412 414
rect 414 412 421 414
rect 408 411 421 412
rect 408 410 418 411
rect 416 409 418 410
rect 420 409 421 411
rect 392 397 393 399
rect 395 397 396 399
rect 360 387 361 389
rect 363 387 364 389
rect 360 386 364 387
rect 392 392 396 397
rect 394 390 396 392
rect 392 385 396 390
rect 394 383 396 385
rect 383 379 396 383
rect 392 378 396 379
rect 400 398 405 400
rect 400 396 402 398
rect 404 396 405 398
rect 400 389 405 396
rect 416 402 421 409
rect 456 414 460 419
rect 456 412 457 414
rect 459 412 460 414
rect 400 387 401 389
rect 403 387 405 389
rect 400 384 405 387
rect 400 378 412 384
rect 456 391 460 412
rect 520 422 524 424
rect 519 420 524 422
rect 519 418 520 420
rect 522 418 524 420
rect 519 416 524 418
rect 471 414 484 415
rect 471 412 472 414
rect 474 412 484 414
rect 471 411 484 412
rect 478 406 484 411
rect 478 404 479 406
rect 481 404 484 406
rect 478 402 484 404
rect 504 401 508 408
rect 504 400 506 401
rect 496 399 506 400
rect 496 397 497 399
rect 499 397 508 399
rect 496 394 508 397
rect 444 389 460 391
rect 444 387 446 389
rect 448 387 460 389
rect 444 386 460 387
rect 464 387 477 391
rect 464 386 469 387
rect 520 390 524 416
rect 584 422 588 424
rect 583 420 588 422
rect 583 418 584 420
rect 586 418 588 420
rect 583 416 588 418
rect 535 414 548 415
rect 535 412 536 414
rect 538 412 548 414
rect 535 411 548 412
rect 542 406 548 411
rect 542 404 543 406
rect 545 404 548 406
rect 542 402 548 404
rect 584 414 588 416
rect 568 401 572 408
rect 584 412 585 414
rect 587 412 588 414
rect 568 400 570 401
rect 560 399 570 400
rect 560 398 572 399
rect 560 396 561 398
rect 563 396 572 398
rect 560 394 572 396
rect 520 388 521 390
rect 523 388 524 390
rect 464 384 466 386
rect 468 384 469 386
rect 464 381 469 384
rect 520 383 524 388
rect 511 382 524 383
rect 464 379 465 381
rect 467 379 469 381
rect 511 380 520 382
rect 522 380 524 382
rect 511 379 524 380
rect 528 387 541 391
rect 528 386 533 387
rect 528 384 530 386
rect 532 384 533 386
rect 528 381 533 384
rect 584 383 588 412
rect 648 422 652 424
rect 647 420 652 422
rect 647 418 648 420
rect 650 418 652 420
rect 647 416 652 418
rect 599 414 612 415
rect 599 412 600 414
rect 602 412 612 414
rect 599 411 612 412
rect 606 406 612 411
rect 606 404 607 406
rect 609 404 612 406
rect 606 402 612 404
rect 632 401 636 408
rect 632 400 634 401
rect 624 399 634 400
rect 624 397 636 399
rect 624 395 625 397
rect 627 395 636 397
rect 624 394 636 395
rect 575 382 588 383
rect 528 379 530 381
rect 532 379 533 381
rect 575 380 584 382
rect 586 380 588 382
rect 575 379 588 380
rect 592 387 605 391
rect 592 386 597 387
rect 592 384 594 386
rect 596 384 597 386
rect 592 381 597 384
rect 648 383 652 416
rect 639 382 652 383
rect 592 379 594 381
rect 596 379 597 381
rect 639 380 648 382
rect 650 380 652 382
rect 639 379 652 380
rect 464 378 469 379
rect 528 378 533 379
rect 592 378 597 379
rect 3 372 656 373
rect 3 370 29 372
rect 31 370 102 372
rect 104 370 133 372
rect 135 370 206 372
rect 208 370 246 372
rect 248 370 278 372
rect 280 370 351 372
rect 353 370 391 372
rect 393 370 436 372
rect 438 370 656 372
rect 3 368 252 370
rect 254 368 656 370
rect 3 361 656 368
rect 3 360 252 361
rect 3 358 10 360
rect 12 358 50 360
rect 52 358 123 360
rect 125 358 154 360
rect 156 358 227 360
rect 229 359 252 360
rect 254 360 656 361
rect 254 359 278 360
rect 229 358 278 359
rect 280 358 351 360
rect 353 358 391 360
rect 393 358 436 360
rect 438 358 656 360
rect 3 357 656 358
rect 7 351 11 352
rect 7 347 20 351
rect 7 345 9 347
rect 7 340 11 345
rect 7 338 9 340
rect 7 326 11 338
rect 39 339 43 344
rect 7 324 8 326
rect 10 324 11 326
rect 7 319 11 324
rect 39 337 40 339
rect 42 337 43 339
rect 39 335 43 337
rect 22 333 43 335
rect 22 331 36 333
rect 38 331 43 333
rect 47 343 52 345
rect 47 341 49 343
rect 51 341 52 343
rect 87 346 99 352
rect 47 339 52 341
rect 47 337 48 339
rect 50 337 52 339
rect 47 336 52 337
rect 47 334 49 336
rect 51 334 52 336
rect 47 332 52 334
rect 79 341 83 344
rect 79 339 80 341
rect 82 339 83 341
rect 7 317 12 319
rect 7 315 9 317
rect 11 315 12 317
rect 7 313 12 315
rect 22 326 43 327
rect 22 324 26 326
rect 28 324 40 326
rect 42 324 43 326
rect 22 323 43 324
rect 39 314 43 323
rect 47 312 51 332
rect 79 335 83 339
rect 70 334 83 335
rect 70 332 76 334
rect 78 332 83 334
rect 70 331 83 332
rect 87 341 92 346
rect 87 339 89 341
rect 91 339 92 341
rect 87 334 92 339
rect 87 332 89 334
rect 91 332 92 334
rect 87 330 92 332
rect 62 326 76 327
rect 62 324 66 326
rect 68 324 76 326
rect 62 323 76 324
rect 47 310 49 312
rect 51 310 59 312
rect 47 306 59 310
rect 71 317 76 323
rect 71 315 72 317
rect 74 315 76 317
rect 71 314 76 315
rect 103 321 108 328
rect 131 343 147 344
rect 131 341 133 343
rect 135 341 147 343
rect 131 339 147 341
rect 143 334 147 339
rect 143 332 144 334
rect 146 332 147 334
rect 103 320 105 321
rect 95 319 105 320
rect 107 319 108 321
rect 95 317 108 319
rect 95 315 97 317
rect 99 315 108 317
rect 95 314 108 315
rect 143 311 147 332
rect 123 310 147 311
rect 123 308 125 310
rect 127 308 147 310
rect 123 307 147 308
rect 151 343 156 345
rect 151 341 153 343
rect 155 341 156 343
rect 191 346 203 352
rect 151 336 156 341
rect 151 334 153 336
rect 155 334 156 336
rect 151 332 156 334
rect 183 341 187 344
rect 183 339 184 341
rect 186 339 187 341
rect 151 326 155 332
rect 151 324 152 326
rect 154 324 155 326
rect 151 312 155 324
rect 183 335 187 339
rect 174 334 187 335
rect 174 332 175 334
rect 177 332 180 334
rect 182 332 187 334
rect 174 331 187 332
rect 191 341 196 346
rect 191 339 193 341
rect 195 339 196 341
rect 191 334 196 339
rect 191 332 193 334
rect 195 332 196 334
rect 191 330 196 332
rect 166 326 180 327
rect 166 324 170 326
rect 172 324 180 326
rect 166 323 180 324
rect 151 310 153 312
rect 155 310 163 312
rect 151 306 163 310
rect 175 317 180 323
rect 175 315 176 317
rect 178 315 180 317
rect 175 314 180 315
rect 207 321 212 328
rect 235 343 251 344
rect 235 341 237 343
rect 239 341 251 343
rect 235 339 251 341
rect 207 320 209 321
rect 199 319 209 320
rect 211 319 212 321
rect 199 317 212 319
rect 199 315 201 317
rect 203 315 212 317
rect 199 314 212 315
rect 247 311 251 339
rect 227 310 251 311
rect 227 308 229 310
rect 231 308 251 310
rect 227 307 251 308
rect 256 343 272 344
rect 256 342 268 343
rect 256 340 257 342
rect 259 341 268 342
rect 270 341 272 343
rect 259 340 272 341
rect 256 339 272 340
rect 256 311 260 339
rect 304 346 316 352
rect 311 342 316 346
rect 311 340 312 342
rect 314 340 316 342
rect 295 321 300 328
rect 311 334 316 340
rect 311 332 312 334
rect 314 332 316 334
rect 311 330 316 332
rect 320 342 324 344
rect 320 340 321 342
rect 323 340 324 342
rect 320 335 324 340
rect 392 351 396 352
rect 383 347 396 351
rect 351 343 356 345
rect 320 334 333 335
rect 320 332 325 334
rect 327 332 333 334
rect 320 331 333 332
rect 295 319 296 321
rect 298 320 300 321
rect 298 319 308 320
rect 295 317 308 319
rect 295 315 303 317
rect 305 315 308 317
rect 295 314 308 315
rect 327 326 341 327
rect 327 324 335 326
rect 337 324 341 326
rect 327 323 341 324
rect 351 341 352 343
rect 354 341 356 343
rect 351 336 356 341
rect 351 334 352 336
rect 354 334 356 336
rect 351 332 356 334
rect 327 318 332 323
rect 327 316 329 318
rect 331 316 332 318
rect 327 314 332 316
rect 256 310 280 311
rect 256 308 276 310
rect 278 308 280 310
rect 352 312 356 332
rect 360 342 364 344
rect 360 340 361 342
rect 363 340 364 342
rect 360 335 364 340
rect 360 333 381 335
rect 360 331 365 333
rect 367 331 381 333
rect 360 326 381 327
rect 360 324 375 326
rect 377 324 381 326
rect 360 323 381 324
rect 394 345 396 347
rect 392 340 396 345
rect 394 338 396 340
rect 360 317 364 323
rect 392 333 396 338
rect 392 331 393 333
rect 395 331 396 333
rect 392 319 396 331
rect 400 346 412 352
rect 464 351 469 352
rect 528 351 533 352
rect 592 351 597 352
rect 464 349 465 351
rect 467 349 469 351
rect 400 342 405 346
rect 400 340 401 342
rect 403 340 405 342
rect 400 334 405 340
rect 464 346 469 349
rect 511 350 524 351
rect 511 348 520 350
rect 522 348 524 350
rect 400 332 402 334
rect 404 332 405 334
rect 400 330 405 332
rect 360 315 361 317
rect 363 315 364 317
rect 360 314 364 315
rect 391 317 396 319
rect 391 315 392 317
rect 394 315 396 317
rect 391 313 396 315
rect 416 321 421 328
rect 464 344 466 346
rect 468 344 469 346
rect 511 347 524 348
rect 444 343 460 344
rect 444 341 446 343
rect 448 341 460 343
rect 444 339 460 341
rect 464 343 469 344
rect 464 339 477 343
rect 416 320 418 321
rect 408 319 418 320
rect 420 319 421 321
rect 408 318 421 319
rect 408 316 413 318
rect 415 316 421 318
rect 408 314 421 316
rect 456 318 460 339
rect 456 316 457 318
rect 459 316 460 318
rect 256 307 280 308
rect 344 310 352 312
rect 354 310 356 312
rect 456 311 460 316
rect 344 309 356 310
rect 344 307 353 309
rect 355 307 356 309
rect 344 306 356 307
rect 436 310 460 311
rect 436 308 438 310
rect 440 308 460 310
rect 478 326 484 328
rect 478 324 479 326
rect 481 324 484 326
rect 478 319 484 324
rect 471 318 484 319
rect 471 316 472 318
rect 474 316 484 318
rect 496 333 508 336
rect 496 331 497 333
rect 499 331 508 333
rect 496 330 506 331
rect 504 329 506 330
rect 504 322 508 329
rect 520 342 524 347
rect 520 340 521 342
rect 523 340 524 342
rect 471 315 484 316
rect 520 314 524 340
rect 528 349 530 351
rect 532 349 533 351
rect 528 346 533 349
rect 575 350 588 351
rect 575 348 584 350
rect 586 348 588 350
rect 528 344 530 346
rect 532 344 533 346
rect 575 347 588 348
rect 528 343 533 344
rect 528 339 541 343
rect 519 312 524 314
rect 436 307 460 308
rect 519 310 520 312
rect 522 310 524 312
rect 519 308 524 310
rect 542 326 548 328
rect 542 324 543 326
rect 545 324 548 326
rect 542 319 548 324
rect 535 318 548 319
rect 535 316 536 318
rect 538 316 548 318
rect 560 333 572 336
rect 560 331 561 333
rect 563 331 572 333
rect 560 330 570 331
rect 568 329 570 330
rect 568 322 572 329
rect 584 318 588 347
rect 592 349 594 351
rect 596 349 597 351
rect 592 346 597 349
rect 639 350 652 351
rect 639 348 648 350
rect 650 348 652 350
rect 592 344 594 346
rect 596 344 597 346
rect 639 347 652 348
rect 592 343 597 344
rect 592 339 605 343
rect 535 315 548 316
rect 584 316 585 318
rect 587 316 588 318
rect 584 314 588 316
rect 583 312 588 314
rect 520 306 524 308
rect 583 310 584 312
rect 586 310 588 312
rect 583 308 588 310
rect 606 326 612 328
rect 606 324 607 326
rect 609 324 612 326
rect 606 319 612 324
rect 599 318 612 319
rect 599 316 600 318
rect 602 316 612 318
rect 624 335 636 336
rect 624 333 625 335
rect 627 333 636 335
rect 624 331 636 333
rect 624 330 634 331
rect 632 329 634 330
rect 632 322 636 329
rect 599 315 612 316
rect 648 314 652 347
rect 647 312 652 314
rect 584 306 588 308
rect 647 310 648 312
rect 650 310 652 312
rect 647 308 652 310
rect 648 306 652 308
rect 3 300 656 301
rect 3 298 10 300
rect 12 298 50 300
rect 52 298 60 300
rect 62 298 90 300
rect 92 298 143 300
rect 145 298 154 300
rect 156 298 164 300
rect 166 298 194 300
rect 196 298 247 300
rect 249 298 258 300
rect 260 298 311 300
rect 313 298 341 300
rect 343 298 351 300
rect 353 298 391 300
rect 393 298 403 300
rect 405 298 456 300
rect 458 298 656 300
rect 3 296 4 298
rect 6 296 656 298
rect 3 290 656 296
rect 3 288 4 290
rect 6 288 656 290
rect 3 286 9 288
rect 11 286 62 288
rect 64 286 92 288
rect 94 286 102 288
rect 104 286 113 288
rect 115 286 166 288
rect 168 286 196 288
rect 198 286 206 288
rect 208 286 246 288
rect 248 286 258 288
rect 260 286 311 288
rect 313 286 341 288
rect 343 286 351 288
rect 353 286 391 288
rect 393 286 403 288
rect 405 286 456 288
rect 458 286 656 288
rect 3 285 656 286
rect 7 278 31 279
rect 7 276 27 278
rect 29 276 31 278
rect 7 275 31 276
rect 7 247 11 275
rect 46 271 59 272
rect 46 269 55 271
rect 57 269 59 271
rect 46 267 59 269
rect 46 265 47 267
rect 49 266 59 267
rect 49 265 51 266
rect 7 245 23 247
rect 7 243 19 245
rect 21 243 23 245
rect 7 242 23 243
rect 46 258 51 265
rect 78 271 83 272
rect 78 269 80 271
rect 82 269 83 271
rect 78 263 83 269
rect 95 276 107 280
rect 95 274 103 276
rect 105 274 107 276
rect 78 262 92 263
rect 78 260 86 262
rect 88 260 89 262
rect 91 260 92 262
rect 78 259 92 260
rect 62 254 67 256
rect 62 252 63 254
rect 65 252 67 254
rect 62 247 67 252
rect 62 245 63 247
rect 65 245 67 247
rect 62 240 67 245
rect 71 254 84 255
rect 71 252 76 254
rect 78 252 81 254
rect 83 252 84 254
rect 71 251 84 252
rect 71 247 75 251
rect 103 262 107 274
rect 103 260 104 262
rect 106 260 107 262
rect 103 254 107 260
rect 71 245 72 247
rect 74 245 75 247
rect 71 242 75 245
rect 102 252 107 254
rect 102 250 103 252
rect 105 250 107 252
rect 102 245 107 250
rect 55 234 67 240
rect 102 243 103 245
rect 105 243 107 245
rect 102 241 107 243
rect 111 278 135 279
rect 111 276 131 278
rect 133 276 135 278
rect 111 275 135 276
rect 111 254 115 275
rect 150 271 163 272
rect 150 269 159 271
rect 161 269 163 271
rect 150 267 163 269
rect 150 265 151 267
rect 153 266 163 267
rect 153 265 155 266
rect 111 252 112 254
rect 114 252 115 254
rect 111 247 115 252
rect 111 245 127 247
rect 111 243 123 245
rect 125 243 127 245
rect 111 242 127 243
rect 150 258 155 265
rect 182 271 187 272
rect 182 269 184 271
rect 186 269 187 271
rect 182 263 187 269
rect 199 276 211 280
rect 344 279 356 280
rect 199 274 207 276
rect 209 274 211 276
rect 182 262 196 263
rect 182 260 190 262
rect 192 260 196 262
rect 182 259 196 260
rect 166 254 171 256
rect 166 252 167 254
rect 169 252 171 254
rect 166 247 171 252
rect 166 245 167 247
rect 169 245 171 247
rect 166 240 171 245
rect 175 254 188 255
rect 175 252 180 254
rect 182 252 188 254
rect 175 251 188 252
rect 175 247 179 251
rect 207 254 211 274
rect 256 278 280 279
rect 256 276 276 278
rect 278 276 280 278
rect 256 275 280 276
rect 215 263 219 272
rect 215 262 236 263
rect 215 260 216 262
rect 218 260 230 262
rect 232 260 236 262
rect 215 259 236 260
rect 246 271 251 273
rect 246 269 247 271
rect 249 269 251 271
rect 246 267 251 269
rect 175 245 176 247
rect 178 245 179 247
rect 175 242 179 245
rect 206 252 211 254
rect 206 250 207 252
rect 209 250 211 252
rect 206 249 211 250
rect 206 247 208 249
rect 210 247 211 249
rect 206 245 211 247
rect 159 234 171 240
rect 206 243 207 245
rect 209 243 211 245
rect 206 241 211 243
rect 215 253 220 255
rect 222 253 236 255
rect 215 251 236 253
rect 215 249 219 251
rect 215 247 216 249
rect 218 247 219 249
rect 247 259 251 267
rect 247 257 248 259
rect 250 257 251 259
rect 215 242 219 247
rect 247 248 251 257
rect 249 246 251 248
rect 247 241 251 246
rect 256 247 260 275
rect 295 270 308 272
rect 295 268 303 270
rect 305 268 308 270
rect 295 267 308 268
rect 295 265 296 267
rect 298 266 308 267
rect 298 265 300 266
rect 256 245 272 247
rect 256 243 257 245
rect 259 243 268 245
rect 270 243 272 245
rect 256 242 272 243
rect 295 258 300 265
rect 327 271 332 272
rect 327 269 329 271
rect 331 269 332 271
rect 327 263 332 269
rect 344 277 353 279
rect 355 277 356 279
rect 344 276 356 277
rect 436 278 460 279
rect 344 274 352 276
rect 354 274 356 276
rect 327 262 341 263
rect 327 260 335 262
rect 337 260 341 262
rect 327 259 341 260
rect 311 254 316 256
rect 311 252 312 254
rect 314 252 316 254
rect 249 239 251 241
rect 238 235 251 239
rect 311 245 316 252
rect 311 243 312 245
rect 314 243 316 245
rect 311 240 316 243
rect 320 254 333 255
rect 320 252 325 254
rect 327 252 333 254
rect 320 251 333 252
rect 320 245 324 251
rect 352 254 356 274
rect 436 276 438 278
rect 440 276 460 278
rect 436 275 460 276
rect 360 270 364 272
rect 360 268 361 270
rect 363 268 364 270
rect 360 263 364 268
rect 360 262 381 263
rect 360 260 375 262
rect 377 260 381 262
rect 360 259 381 260
rect 391 271 396 273
rect 391 269 392 271
rect 394 269 396 271
rect 391 267 396 269
rect 320 243 321 245
rect 323 243 324 245
rect 320 242 324 243
rect 351 252 356 254
rect 351 250 352 252
rect 354 250 356 252
rect 351 245 356 250
rect 247 234 251 235
rect 304 234 316 240
rect 351 243 352 245
rect 354 243 356 245
rect 351 241 356 243
rect 360 253 365 255
rect 367 253 381 255
rect 360 251 381 253
rect 360 245 364 251
rect 392 255 396 267
rect 408 271 421 272
rect 408 269 412 271
rect 414 269 421 271
rect 408 267 421 269
rect 408 266 418 267
rect 416 265 418 266
rect 420 265 421 267
rect 392 253 393 255
rect 395 253 396 255
rect 360 243 361 245
rect 363 243 364 245
rect 360 242 364 243
rect 392 248 396 253
rect 394 246 396 248
rect 392 241 396 246
rect 394 239 396 241
rect 383 235 396 239
rect 392 234 396 235
rect 400 254 405 256
rect 400 252 402 254
rect 404 252 405 254
rect 400 245 405 252
rect 416 258 421 265
rect 456 270 460 275
rect 456 268 457 270
rect 459 268 460 270
rect 400 243 401 245
rect 403 243 405 245
rect 400 240 405 243
rect 400 234 412 240
rect 456 247 460 268
rect 520 278 524 280
rect 519 276 524 278
rect 519 274 520 276
rect 522 274 524 276
rect 519 272 524 274
rect 471 270 484 271
rect 471 268 472 270
rect 474 268 484 270
rect 471 267 484 268
rect 478 262 484 267
rect 478 260 479 262
rect 481 260 484 262
rect 478 258 484 260
rect 504 257 508 264
rect 504 256 506 257
rect 496 255 506 256
rect 496 253 497 255
rect 499 253 508 255
rect 496 250 508 253
rect 444 245 460 247
rect 444 243 446 245
rect 448 243 460 245
rect 444 242 460 243
rect 464 243 477 247
rect 464 242 469 243
rect 520 246 524 272
rect 584 278 588 280
rect 583 276 588 278
rect 583 274 584 276
rect 586 274 588 276
rect 583 272 588 274
rect 535 270 548 271
rect 535 268 536 270
rect 538 268 548 270
rect 535 267 548 268
rect 542 262 548 267
rect 542 260 543 262
rect 545 260 548 262
rect 542 258 548 260
rect 584 270 588 272
rect 568 257 572 264
rect 584 268 585 270
rect 587 268 588 270
rect 568 256 570 257
rect 560 255 570 256
rect 560 253 561 255
rect 563 253 572 255
rect 560 250 572 253
rect 520 244 521 246
rect 523 244 524 246
rect 464 240 466 242
rect 468 240 469 242
rect 464 237 469 240
rect 520 239 524 244
rect 511 238 524 239
rect 464 235 465 237
rect 467 235 469 237
rect 511 236 520 238
rect 522 236 524 238
rect 511 235 524 236
rect 528 243 541 247
rect 528 242 533 243
rect 528 240 530 242
rect 532 240 533 242
rect 528 237 533 240
rect 584 239 588 268
rect 648 278 652 280
rect 647 276 652 278
rect 647 274 648 276
rect 650 274 652 276
rect 647 272 652 274
rect 599 270 612 271
rect 599 268 600 270
rect 602 268 612 270
rect 599 267 612 268
rect 606 262 612 267
rect 606 260 607 262
rect 609 260 612 262
rect 606 258 612 260
rect 632 257 636 264
rect 632 256 634 257
rect 624 255 634 256
rect 624 253 636 255
rect 624 251 625 253
rect 627 251 636 253
rect 624 250 636 251
rect 575 238 588 239
rect 528 235 529 237
rect 531 235 533 237
rect 575 236 584 238
rect 586 236 588 238
rect 575 235 588 236
rect 592 243 605 247
rect 592 242 597 243
rect 592 240 594 242
rect 596 240 597 242
rect 592 237 597 240
rect 648 239 652 272
rect 639 238 652 239
rect 592 235 594 237
rect 596 235 597 237
rect 639 236 648 238
rect 650 236 652 238
rect 639 235 652 236
rect 464 234 469 235
rect 528 234 533 235
rect 592 234 597 235
rect 3 228 656 229
rect 3 226 29 228
rect 31 226 102 228
rect 104 226 133 228
rect 135 226 206 228
rect 208 226 246 228
rect 248 227 278 228
rect 248 226 252 227
rect 3 225 252 226
rect 254 226 278 227
rect 280 226 351 228
rect 353 226 391 228
rect 393 226 436 228
rect 438 226 656 228
rect 254 225 656 226
rect 3 217 656 225
rect 3 216 252 217
rect 3 214 10 216
rect 12 214 50 216
rect 52 214 123 216
rect 125 214 154 216
rect 156 214 227 216
rect 229 215 252 216
rect 254 216 656 217
rect 254 215 278 216
rect 229 214 278 215
rect 280 214 351 216
rect 353 214 391 216
rect 393 214 436 216
rect 438 214 656 216
rect 3 213 656 214
rect 7 207 11 208
rect 7 203 20 207
rect 7 201 9 203
rect 7 196 11 201
rect 7 194 9 196
rect 7 184 11 194
rect 39 195 43 200
rect 7 182 8 184
rect 10 182 11 184
rect 7 175 11 182
rect 39 193 40 195
rect 42 193 43 195
rect 39 191 43 193
rect 22 189 43 191
rect 22 187 36 189
rect 38 187 43 189
rect 47 199 52 201
rect 47 197 49 199
rect 51 197 52 199
rect 87 202 99 208
rect 47 195 52 197
rect 47 193 48 195
rect 50 193 52 195
rect 47 192 52 193
rect 47 190 49 192
rect 51 190 52 192
rect 47 188 52 190
rect 79 197 83 200
rect 79 195 80 197
rect 82 195 83 197
rect 7 173 12 175
rect 7 171 9 173
rect 11 171 12 173
rect 7 169 12 171
rect 22 182 43 183
rect 22 180 26 182
rect 28 180 40 182
rect 42 180 43 182
rect 22 179 43 180
rect 39 170 43 179
rect 47 168 51 188
rect 79 191 83 195
rect 70 190 83 191
rect 70 188 76 190
rect 78 188 83 190
rect 70 187 83 188
rect 87 197 92 202
rect 87 195 89 197
rect 91 195 92 197
rect 87 190 92 195
rect 87 188 89 190
rect 91 188 92 190
rect 87 186 92 188
rect 62 182 76 183
rect 62 180 66 182
rect 68 180 76 182
rect 62 179 76 180
rect 47 166 49 168
rect 51 166 59 168
rect 47 162 59 166
rect 71 173 76 179
rect 71 171 72 173
rect 74 171 76 173
rect 71 170 76 171
rect 103 177 108 184
rect 131 199 147 200
rect 131 197 133 199
rect 135 197 147 199
rect 131 195 147 197
rect 143 190 147 195
rect 143 188 144 190
rect 146 188 147 190
rect 103 176 105 177
rect 95 175 105 176
rect 107 175 108 177
rect 95 173 108 175
rect 95 171 97 173
rect 99 171 108 173
rect 95 170 108 171
rect 143 167 147 188
rect 123 166 147 167
rect 123 164 125 166
rect 127 164 147 166
rect 123 163 147 164
rect 151 199 156 201
rect 151 197 153 199
rect 155 197 156 199
rect 191 202 203 208
rect 151 192 156 197
rect 151 190 153 192
rect 155 190 156 192
rect 151 188 156 190
rect 183 197 187 200
rect 183 195 184 197
rect 186 195 187 197
rect 151 182 155 188
rect 151 180 152 182
rect 154 180 155 182
rect 151 168 155 180
rect 183 191 187 195
rect 174 190 187 191
rect 174 188 175 190
rect 177 188 180 190
rect 182 188 187 190
rect 174 187 187 188
rect 191 197 196 202
rect 191 195 193 197
rect 195 195 196 197
rect 191 190 196 195
rect 191 188 193 190
rect 195 188 196 190
rect 191 186 196 188
rect 166 182 180 183
rect 166 180 170 182
rect 172 180 177 182
rect 179 180 180 182
rect 166 179 180 180
rect 151 166 153 168
rect 155 166 163 168
rect 151 162 163 166
rect 175 173 180 179
rect 175 171 176 173
rect 178 171 180 173
rect 175 170 180 171
rect 207 177 212 184
rect 235 199 251 200
rect 235 197 237 199
rect 239 198 251 199
rect 239 197 243 198
rect 235 196 243 197
rect 245 196 251 198
rect 235 195 251 196
rect 207 176 209 177
rect 199 175 209 176
rect 211 175 212 177
rect 199 173 212 175
rect 199 171 201 173
rect 203 171 212 173
rect 199 170 212 171
rect 247 167 251 195
rect 227 166 251 167
rect 227 164 229 166
rect 231 164 251 166
rect 227 163 251 164
rect 256 199 272 200
rect 256 198 268 199
rect 256 196 257 198
rect 259 197 268 198
rect 270 197 272 199
rect 259 196 272 197
rect 256 195 272 196
rect 256 167 260 195
rect 304 202 316 208
rect 311 198 316 202
rect 311 196 312 198
rect 314 196 316 198
rect 295 177 300 184
rect 311 190 316 196
rect 311 188 312 190
rect 314 188 316 190
rect 311 186 316 188
rect 320 198 324 200
rect 320 196 321 198
rect 323 196 324 198
rect 320 191 324 196
rect 392 207 396 208
rect 383 203 396 207
rect 351 199 356 201
rect 320 190 333 191
rect 320 188 325 190
rect 327 188 333 190
rect 320 187 333 188
rect 295 175 296 177
rect 298 176 300 177
rect 298 175 308 176
rect 295 174 308 175
rect 295 172 303 174
rect 305 172 308 174
rect 295 170 308 172
rect 327 182 341 183
rect 327 180 335 182
rect 337 180 341 182
rect 327 179 341 180
rect 351 197 352 199
rect 354 197 356 199
rect 351 192 356 197
rect 351 190 352 192
rect 354 190 356 192
rect 351 188 356 190
rect 327 173 332 179
rect 327 171 329 173
rect 331 171 332 173
rect 327 170 332 171
rect 256 166 280 167
rect 256 164 276 166
rect 278 164 280 166
rect 352 168 356 188
rect 360 198 364 200
rect 360 196 361 198
rect 363 196 364 198
rect 360 191 364 196
rect 360 189 381 191
rect 360 187 365 189
rect 367 187 381 189
rect 360 182 381 183
rect 360 180 375 182
rect 377 180 381 182
rect 360 179 381 180
rect 394 201 396 203
rect 392 196 396 201
rect 394 194 396 196
rect 360 173 364 179
rect 392 189 396 194
rect 392 187 393 189
rect 395 187 396 189
rect 392 175 396 187
rect 400 202 412 208
rect 464 207 469 208
rect 528 207 533 208
rect 592 207 597 208
rect 464 205 465 207
rect 467 205 469 207
rect 400 198 405 202
rect 400 196 401 198
rect 403 196 405 198
rect 400 190 405 196
rect 464 202 469 205
rect 511 206 524 207
rect 511 204 520 206
rect 522 204 524 206
rect 400 188 402 190
rect 404 188 405 190
rect 400 186 405 188
rect 360 171 361 173
rect 363 171 364 173
rect 360 170 364 171
rect 391 173 396 175
rect 391 171 392 173
rect 394 171 396 173
rect 391 169 396 171
rect 416 177 421 184
rect 464 200 466 202
rect 468 200 469 202
rect 511 203 524 204
rect 444 199 460 200
rect 444 197 446 199
rect 448 197 460 199
rect 444 195 460 197
rect 464 199 469 200
rect 464 195 477 199
rect 416 176 418 177
rect 408 175 418 176
rect 420 175 421 177
rect 408 174 421 175
rect 408 172 412 174
rect 414 172 421 174
rect 408 170 421 172
rect 456 174 460 195
rect 456 172 457 174
rect 459 172 460 174
rect 256 163 280 164
rect 344 166 352 168
rect 354 166 356 168
rect 456 167 460 172
rect 344 165 356 166
rect 344 163 353 165
rect 355 163 356 165
rect 344 162 356 163
rect 436 166 460 167
rect 436 164 438 166
rect 440 164 460 166
rect 478 182 484 184
rect 478 180 479 182
rect 481 180 484 182
rect 478 175 484 180
rect 471 174 484 175
rect 471 172 472 174
rect 474 172 484 174
rect 496 189 508 192
rect 496 187 497 189
rect 499 187 508 189
rect 496 186 506 187
rect 504 185 506 186
rect 504 178 508 185
rect 520 198 524 203
rect 520 196 521 198
rect 523 196 524 198
rect 471 171 484 172
rect 520 170 524 196
rect 528 205 529 207
rect 531 205 533 207
rect 528 202 533 205
rect 575 206 588 207
rect 575 204 584 206
rect 586 204 588 206
rect 528 200 530 202
rect 532 200 533 202
rect 575 203 588 204
rect 528 199 533 200
rect 528 195 541 199
rect 519 168 524 170
rect 436 163 460 164
rect 519 166 520 168
rect 522 166 524 168
rect 519 164 524 166
rect 542 182 548 184
rect 542 180 543 182
rect 545 180 548 182
rect 542 175 548 180
rect 535 174 548 175
rect 535 172 536 174
rect 538 172 548 174
rect 560 189 572 192
rect 560 187 561 189
rect 563 187 572 189
rect 560 186 570 187
rect 568 185 570 186
rect 568 178 572 185
rect 584 174 588 203
rect 592 205 594 207
rect 596 205 597 207
rect 592 202 597 205
rect 639 206 652 207
rect 639 204 648 206
rect 650 204 652 206
rect 592 200 594 202
rect 596 200 597 202
rect 639 203 652 204
rect 592 199 597 200
rect 592 195 605 199
rect 535 171 548 172
rect 584 172 585 174
rect 587 172 588 174
rect 584 170 588 172
rect 583 168 588 170
rect 520 162 524 164
rect 583 166 584 168
rect 586 166 588 168
rect 583 164 588 166
rect 606 182 612 184
rect 606 180 607 182
rect 609 180 612 182
rect 606 175 612 180
rect 599 174 612 175
rect 599 172 600 174
rect 602 172 612 174
rect 624 191 636 192
rect 624 189 625 191
rect 627 189 636 191
rect 624 187 636 189
rect 624 186 634 187
rect 632 185 634 186
rect 632 178 636 185
rect 599 171 612 172
rect 648 170 652 203
rect 647 168 652 170
rect 584 162 588 164
rect 647 166 648 168
rect 650 166 652 168
rect 647 164 652 166
rect 648 162 652 164
rect 3 156 656 157
rect 3 154 4 156
rect 6 154 10 156
rect 12 154 50 156
rect 52 154 60 156
rect 62 154 90 156
rect 92 154 143 156
rect 145 154 154 156
rect 156 154 164 156
rect 166 154 194 156
rect 196 154 247 156
rect 249 154 258 156
rect 260 154 311 156
rect 313 154 341 156
rect 343 154 351 156
rect 353 154 391 156
rect 393 154 403 156
rect 405 154 456 156
rect 458 154 656 156
rect 3 146 656 154
rect 3 144 4 146
rect 6 144 656 146
rect 3 142 9 144
rect 11 142 62 144
rect 64 142 92 144
rect 94 142 102 144
rect 104 142 113 144
rect 115 142 166 144
rect 168 142 196 144
rect 198 142 206 144
rect 208 142 246 144
rect 248 142 258 144
rect 260 142 311 144
rect 313 142 341 144
rect 343 142 351 144
rect 353 142 391 144
rect 393 142 403 144
rect 405 142 456 144
rect 458 142 656 144
rect 3 141 656 142
rect 7 134 31 135
rect 7 132 27 134
rect 29 132 31 134
rect 7 131 31 132
rect 7 103 11 131
rect 46 127 59 128
rect 46 125 55 127
rect 57 125 59 127
rect 46 123 59 125
rect 46 121 47 123
rect 49 122 59 123
rect 49 121 51 122
rect 7 101 23 103
rect 7 99 19 101
rect 21 99 23 101
rect 7 98 23 99
rect 46 114 51 121
rect 78 127 83 128
rect 78 125 80 127
rect 82 125 83 127
rect 78 119 83 125
rect 95 132 107 136
rect 95 130 103 132
rect 105 130 107 132
rect 78 118 92 119
rect 78 116 81 118
rect 83 116 86 118
rect 88 116 92 118
rect 78 115 92 116
rect 62 110 67 112
rect 62 108 63 110
rect 65 108 67 110
rect 62 103 67 108
rect 62 101 63 103
rect 65 101 67 103
rect 62 96 67 101
rect 71 110 84 111
rect 71 108 76 110
rect 78 108 81 110
rect 83 108 84 110
rect 71 107 84 108
rect 71 103 75 107
rect 103 118 107 130
rect 103 116 104 118
rect 106 116 107 118
rect 103 110 107 116
rect 71 101 72 103
rect 74 101 75 103
rect 71 98 75 101
rect 102 108 107 110
rect 102 106 103 108
rect 105 106 107 108
rect 102 101 107 106
rect 55 90 67 96
rect 102 99 103 101
rect 105 99 107 101
rect 102 97 107 99
rect 111 134 135 135
rect 111 132 131 134
rect 133 132 135 134
rect 111 131 135 132
rect 111 110 115 131
rect 150 127 163 128
rect 150 125 159 127
rect 161 125 163 127
rect 150 123 163 125
rect 150 121 151 123
rect 153 122 163 123
rect 153 121 155 122
rect 111 108 112 110
rect 114 108 115 110
rect 111 103 115 108
rect 111 101 127 103
rect 111 99 123 101
rect 125 99 127 101
rect 111 98 127 99
rect 150 114 155 121
rect 182 127 187 128
rect 182 125 184 127
rect 186 125 187 127
rect 182 119 187 125
rect 199 132 211 136
rect 344 135 356 136
rect 199 130 207 132
rect 209 130 211 132
rect 182 118 196 119
rect 182 116 190 118
rect 192 116 196 118
rect 182 115 196 116
rect 166 110 171 112
rect 166 108 167 110
rect 169 108 171 110
rect 166 103 171 108
rect 166 101 167 103
rect 169 101 171 103
rect 166 96 171 101
rect 175 110 188 111
rect 175 108 180 110
rect 182 108 188 110
rect 175 107 188 108
rect 175 103 179 107
rect 207 110 211 130
rect 256 134 280 135
rect 256 132 276 134
rect 278 132 280 134
rect 256 131 280 132
rect 215 119 219 128
rect 215 118 236 119
rect 215 116 216 118
rect 218 116 230 118
rect 232 116 236 118
rect 215 115 236 116
rect 246 127 251 129
rect 246 125 247 127
rect 249 125 251 127
rect 246 123 251 125
rect 175 101 176 103
rect 178 101 179 103
rect 175 98 179 101
rect 206 108 211 110
rect 206 106 207 108
rect 209 106 211 108
rect 206 105 211 106
rect 206 103 208 105
rect 210 103 211 105
rect 206 101 211 103
rect 159 90 171 96
rect 206 99 207 101
rect 209 99 211 101
rect 206 97 211 99
rect 215 109 220 111
rect 222 109 236 111
rect 215 107 236 109
rect 215 105 219 107
rect 215 103 216 105
rect 218 103 219 105
rect 247 120 251 123
rect 247 118 248 120
rect 250 118 251 120
rect 215 98 219 103
rect 247 104 251 118
rect 249 102 251 104
rect 247 97 251 102
rect 256 103 260 131
rect 295 126 308 128
rect 295 124 303 126
rect 305 124 308 126
rect 295 123 308 124
rect 295 121 296 123
rect 298 122 308 123
rect 298 121 300 122
rect 256 101 272 103
rect 256 99 257 101
rect 259 99 268 101
rect 270 99 272 101
rect 256 98 272 99
rect 295 114 300 121
rect 327 126 332 128
rect 327 124 329 126
rect 331 124 332 126
rect 327 119 332 124
rect 344 133 353 135
rect 355 133 356 135
rect 344 132 356 133
rect 436 134 460 135
rect 344 130 352 132
rect 354 130 356 132
rect 327 118 341 119
rect 327 116 335 118
rect 337 116 341 118
rect 327 115 341 116
rect 311 110 316 112
rect 311 108 312 110
rect 314 108 316 110
rect 249 95 251 97
rect 238 91 251 95
rect 311 101 316 108
rect 311 99 312 101
rect 314 99 316 101
rect 311 96 316 99
rect 320 110 333 111
rect 320 108 325 110
rect 327 108 333 110
rect 320 107 333 108
rect 320 101 324 107
rect 352 110 356 130
rect 436 132 438 134
rect 440 132 460 134
rect 436 131 460 132
rect 360 127 364 128
rect 360 125 361 127
rect 363 125 364 127
rect 360 119 364 125
rect 360 118 381 119
rect 360 116 375 118
rect 377 116 381 118
rect 360 115 381 116
rect 391 127 396 129
rect 391 125 392 127
rect 394 125 396 127
rect 391 123 396 125
rect 320 99 321 101
rect 323 99 324 101
rect 320 98 324 99
rect 351 108 356 110
rect 351 106 352 108
rect 354 106 356 108
rect 351 101 356 106
rect 247 90 251 91
rect 304 90 316 96
rect 351 99 352 101
rect 354 99 356 101
rect 351 97 356 99
rect 360 109 365 111
rect 367 109 381 111
rect 360 107 381 109
rect 360 101 364 107
rect 392 110 396 123
rect 408 127 421 128
rect 408 125 412 127
rect 414 125 421 127
rect 408 123 421 125
rect 408 122 418 123
rect 416 121 418 122
rect 420 121 421 123
rect 392 108 393 110
rect 395 108 396 110
rect 360 99 361 101
rect 363 99 364 101
rect 360 98 364 99
rect 392 104 396 108
rect 394 102 396 104
rect 392 97 396 102
rect 394 95 396 97
rect 383 91 396 95
rect 392 90 396 91
rect 400 110 405 112
rect 400 108 402 110
rect 404 108 405 110
rect 400 101 405 108
rect 416 114 421 121
rect 456 126 460 131
rect 456 124 457 126
rect 459 124 460 126
rect 400 99 401 101
rect 403 99 405 101
rect 400 96 405 99
rect 400 90 412 96
rect 456 103 460 124
rect 520 134 524 136
rect 519 132 524 134
rect 519 130 520 132
rect 522 130 524 132
rect 519 128 524 130
rect 471 126 484 127
rect 471 124 472 126
rect 474 124 484 126
rect 471 123 484 124
rect 478 118 484 123
rect 478 116 479 118
rect 481 116 484 118
rect 478 114 484 116
rect 504 113 508 120
rect 504 112 506 113
rect 496 111 506 112
rect 496 110 508 111
rect 496 108 497 110
rect 499 108 508 110
rect 496 106 508 108
rect 444 101 460 103
rect 444 99 446 101
rect 448 99 460 101
rect 444 98 460 99
rect 464 99 477 103
rect 464 98 469 99
rect 520 102 524 128
rect 584 134 588 136
rect 583 132 588 134
rect 583 130 584 132
rect 586 130 588 132
rect 583 128 588 130
rect 535 126 548 127
rect 535 124 536 126
rect 538 124 548 126
rect 535 123 548 124
rect 542 118 548 123
rect 542 116 543 118
rect 545 116 548 118
rect 542 114 548 116
rect 584 126 588 128
rect 568 113 572 120
rect 584 124 585 126
rect 587 124 588 126
rect 568 112 570 113
rect 560 111 570 112
rect 560 110 572 111
rect 560 108 561 110
rect 563 108 572 110
rect 560 106 572 108
rect 520 100 521 102
rect 523 100 524 102
rect 464 96 466 98
rect 468 96 469 98
rect 464 93 469 96
rect 520 95 524 100
rect 511 94 524 95
rect 464 91 465 93
rect 467 91 469 93
rect 511 92 520 94
rect 522 92 524 94
rect 511 91 524 92
rect 528 99 541 103
rect 528 98 533 99
rect 528 96 530 98
rect 532 96 533 98
rect 528 93 533 96
rect 584 95 588 124
rect 648 134 652 136
rect 647 132 652 134
rect 647 130 648 132
rect 650 130 652 132
rect 647 128 652 130
rect 599 126 612 127
rect 599 124 600 126
rect 602 124 612 126
rect 599 123 612 124
rect 606 118 612 123
rect 606 116 607 118
rect 609 116 612 118
rect 606 114 612 116
rect 632 113 636 120
rect 632 112 634 113
rect 624 111 634 112
rect 624 109 636 111
rect 624 107 625 109
rect 627 107 636 109
rect 624 106 636 107
rect 575 94 588 95
rect 528 91 529 93
rect 531 91 533 93
rect 575 92 584 94
rect 586 92 588 94
rect 575 91 588 92
rect 592 99 605 103
rect 592 98 597 99
rect 592 96 594 98
rect 596 96 597 98
rect 592 93 597 96
rect 648 95 652 128
rect 639 94 652 95
rect 592 91 594 93
rect 596 91 597 93
rect 639 92 648 94
rect 650 92 652 94
rect 639 91 652 92
rect 464 90 469 91
rect 528 90 533 91
rect 592 90 597 91
rect 3 84 656 85
rect 3 82 29 84
rect 31 82 102 84
rect 104 82 133 84
rect 135 82 206 84
rect 208 82 246 84
rect 248 82 278 84
rect 280 82 351 84
rect 353 82 391 84
rect 393 82 436 84
rect 438 82 656 84
rect 3 80 252 82
rect 254 80 656 82
rect 3 72 656 80
rect 3 70 10 72
rect 12 70 50 72
rect 52 70 123 72
rect 125 70 154 72
rect 156 70 227 72
rect 229 70 278 72
rect 280 70 351 72
rect 353 70 391 72
rect 393 70 436 72
rect 438 70 656 72
rect 3 69 656 70
rect 7 63 11 64
rect 7 59 20 63
rect 7 57 9 59
rect 7 52 11 57
rect 7 50 9 52
rect 7 38 11 50
rect 39 51 43 56
rect 7 36 8 38
rect 10 36 11 38
rect 7 31 11 36
rect 39 49 40 51
rect 42 49 43 51
rect 39 47 43 49
rect 22 45 43 47
rect 22 43 36 45
rect 38 43 43 45
rect 47 55 52 57
rect 47 53 49 55
rect 51 53 52 55
rect 87 58 99 64
rect 47 51 52 53
rect 47 49 48 51
rect 50 49 52 51
rect 47 48 52 49
rect 47 46 49 48
rect 51 46 52 48
rect 47 44 52 46
rect 79 53 83 56
rect 79 51 80 53
rect 82 51 83 53
rect 7 29 12 31
rect 7 27 9 29
rect 11 27 12 29
rect 7 25 12 27
rect 22 38 43 39
rect 22 36 26 38
rect 28 36 40 38
rect 42 36 43 38
rect 22 35 43 36
rect 39 26 43 35
rect 47 24 51 44
rect 79 47 83 51
rect 70 46 83 47
rect 70 44 76 46
rect 78 44 83 46
rect 70 43 83 44
rect 87 53 92 58
rect 87 51 89 53
rect 91 51 92 53
rect 87 46 92 51
rect 87 44 89 46
rect 91 44 92 46
rect 87 42 92 44
rect 62 38 76 39
rect 62 36 66 38
rect 68 36 76 38
rect 62 35 76 36
rect 47 22 49 24
rect 51 22 59 24
rect 47 18 59 22
rect 71 29 76 35
rect 71 27 72 29
rect 74 27 76 29
rect 71 26 76 27
rect 103 33 108 40
rect 131 55 147 56
rect 131 53 133 55
rect 135 53 147 55
rect 131 51 147 53
rect 143 46 147 51
rect 143 44 144 46
rect 146 44 147 46
rect 103 32 105 33
rect 95 31 105 32
rect 107 31 108 33
rect 95 29 108 31
rect 95 27 97 29
rect 99 27 108 29
rect 95 26 108 27
rect 143 23 147 44
rect 123 22 147 23
rect 123 20 125 22
rect 127 20 147 22
rect 123 19 147 20
rect 151 55 156 57
rect 151 53 153 55
rect 155 53 156 55
rect 191 58 203 64
rect 151 48 156 53
rect 151 46 153 48
rect 155 46 156 48
rect 151 44 156 46
rect 183 53 187 56
rect 183 51 184 53
rect 186 51 187 53
rect 151 38 155 44
rect 151 36 152 38
rect 154 36 155 38
rect 151 24 155 36
rect 183 47 187 51
rect 174 46 187 47
rect 174 44 175 46
rect 177 44 180 46
rect 182 44 187 46
rect 174 43 187 44
rect 191 53 196 58
rect 191 51 193 53
rect 195 51 196 53
rect 191 46 196 51
rect 191 44 193 46
rect 195 44 196 46
rect 191 42 196 44
rect 166 38 180 39
rect 166 36 170 38
rect 172 36 180 38
rect 166 35 180 36
rect 151 22 153 24
rect 155 22 163 24
rect 151 18 163 22
rect 175 29 180 35
rect 175 27 176 29
rect 178 27 180 29
rect 175 26 180 27
rect 207 33 212 40
rect 235 55 251 56
rect 235 53 237 55
rect 239 53 251 55
rect 235 51 251 53
rect 247 45 251 51
rect 247 43 248 45
rect 250 43 251 45
rect 207 32 209 33
rect 199 31 209 32
rect 211 31 212 33
rect 199 29 212 31
rect 199 27 201 29
rect 203 27 212 29
rect 199 26 212 27
rect 247 23 251 43
rect 227 22 251 23
rect 227 20 229 22
rect 231 20 251 22
rect 227 19 251 20
rect 256 55 272 56
rect 256 54 268 55
rect 256 52 257 54
rect 259 53 268 54
rect 270 53 272 55
rect 259 52 272 53
rect 256 51 272 52
rect 256 23 260 51
rect 304 58 316 64
rect 311 54 316 58
rect 311 52 312 54
rect 314 52 316 54
rect 295 33 300 40
rect 311 46 316 52
rect 311 44 312 46
rect 314 44 316 46
rect 311 42 316 44
rect 320 54 324 56
rect 320 52 321 54
rect 323 52 324 54
rect 320 47 324 52
rect 392 63 396 64
rect 383 59 396 63
rect 351 55 356 57
rect 320 46 333 47
rect 320 44 325 46
rect 327 44 333 46
rect 320 43 333 44
rect 295 31 296 33
rect 298 32 300 33
rect 298 31 308 32
rect 295 29 308 31
rect 295 27 303 29
rect 305 27 308 29
rect 295 26 308 27
rect 327 38 341 39
rect 327 36 335 38
rect 337 36 341 38
rect 327 35 341 36
rect 351 53 352 55
rect 354 53 356 55
rect 351 48 356 53
rect 351 46 352 48
rect 354 46 356 48
rect 351 44 356 46
rect 327 29 332 35
rect 327 27 329 29
rect 331 27 332 29
rect 327 26 332 27
rect 256 22 280 23
rect 256 20 276 22
rect 278 20 280 22
rect 352 24 356 44
rect 360 55 364 56
rect 360 53 361 55
rect 363 53 364 55
rect 360 47 364 53
rect 360 45 381 47
rect 360 43 365 45
rect 367 43 381 45
rect 360 38 381 39
rect 360 36 375 38
rect 377 36 381 38
rect 360 35 381 36
rect 394 57 396 59
rect 392 52 396 57
rect 394 50 396 52
rect 360 29 364 35
rect 392 45 396 50
rect 392 43 393 45
rect 395 43 396 45
rect 392 31 396 43
rect 400 58 412 64
rect 464 63 469 64
rect 528 63 533 64
rect 592 63 597 64
rect 464 61 465 63
rect 467 61 469 63
rect 400 54 405 58
rect 400 52 401 54
rect 403 52 405 54
rect 400 46 405 52
rect 464 58 469 61
rect 511 62 524 63
rect 511 60 520 62
rect 522 60 524 62
rect 400 44 402 46
rect 404 44 405 46
rect 400 42 405 44
rect 360 27 361 29
rect 363 27 364 29
rect 360 26 364 27
rect 391 29 396 31
rect 391 27 392 29
rect 394 27 396 29
rect 391 25 396 27
rect 416 33 421 40
rect 464 56 466 58
rect 468 56 469 58
rect 511 59 524 60
rect 444 55 460 56
rect 444 53 446 55
rect 448 53 460 55
rect 444 51 460 53
rect 464 55 469 56
rect 464 51 477 55
rect 416 32 418 33
rect 408 31 418 32
rect 420 31 421 33
rect 408 30 421 31
rect 408 28 412 30
rect 414 28 421 30
rect 408 26 421 28
rect 456 30 460 51
rect 456 28 457 30
rect 459 28 460 30
rect 256 19 280 20
rect 344 22 352 24
rect 354 22 356 24
rect 456 23 460 28
rect 344 21 356 22
rect 344 19 353 21
rect 355 19 356 21
rect 344 18 356 19
rect 436 22 460 23
rect 436 20 438 22
rect 440 20 460 22
rect 478 38 484 40
rect 478 36 479 38
rect 481 36 484 38
rect 478 31 484 36
rect 471 30 484 31
rect 471 28 478 30
rect 480 28 484 30
rect 496 45 508 48
rect 496 43 497 45
rect 499 43 508 45
rect 496 42 506 43
rect 504 41 506 42
rect 504 34 508 41
rect 520 54 524 59
rect 520 52 521 54
rect 523 52 524 54
rect 471 27 484 28
rect 520 26 524 52
rect 528 61 530 63
rect 532 61 533 63
rect 528 58 533 61
rect 575 62 588 63
rect 575 60 584 62
rect 586 60 588 62
rect 528 56 530 58
rect 532 56 533 58
rect 575 59 588 60
rect 528 55 533 56
rect 528 51 541 55
rect 519 24 524 26
rect 436 19 460 20
rect 519 22 520 24
rect 522 22 524 24
rect 519 20 524 22
rect 542 38 548 40
rect 542 36 543 38
rect 545 36 548 38
rect 542 31 548 36
rect 535 30 548 31
rect 535 28 536 30
rect 538 28 548 30
rect 560 45 572 48
rect 560 43 561 45
rect 563 43 572 45
rect 560 42 570 43
rect 568 41 570 42
rect 568 34 572 41
rect 584 30 588 59
rect 592 61 594 63
rect 596 61 597 63
rect 592 58 597 61
rect 639 62 652 63
rect 639 60 648 62
rect 650 60 652 62
rect 592 56 594 58
rect 596 56 597 58
rect 639 59 652 60
rect 592 55 597 56
rect 592 51 605 55
rect 535 27 548 28
rect 584 28 585 30
rect 587 28 588 30
rect 584 26 588 28
rect 583 24 588 26
rect 520 18 524 20
rect 583 22 584 24
rect 586 22 588 24
rect 583 20 588 22
rect 606 38 612 40
rect 606 36 607 38
rect 609 36 612 38
rect 606 31 612 36
rect 599 30 612 31
rect 599 28 600 30
rect 602 28 612 30
rect 624 47 636 48
rect 624 45 625 47
rect 627 45 636 47
rect 624 43 636 45
rect 624 42 634 43
rect 632 41 634 42
rect 632 34 636 41
rect 599 27 612 28
rect 648 26 652 59
rect 647 24 652 26
rect 584 18 588 20
rect 647 22 648 24
rect 650 22 652 24
rect 647 20 652 22
rect 648 18 652 20
rect 3 12 656 13
rect 3 10 10 12
rect 12 10 50 12
rect 52 10 60 12
rect 62 10 90 12
rect 92 10 143 12
rect 145 10 154 12
rect 156 10 164 12
rect 166 10 194 12
rect 196 10 247 12
rect 249 10 258 12
rect 260 10 311 12
rect 313 10 341 12
rect 343 10 351 12
rect 353 10 391 12
rect 393 10 403 12
rect 405 10 456 12
rect 458 10 656 12
rect 3 8 4 10
rect 6 8 656 10
rect 3 5 656 8
<< alu2 >>
rect 3 578 7 579
rect 3 576 4 578
rect 6 576 7 578
rect 3 575 7 576
rect 352 567 539 568
rect 352 565 353 567
rect 355 565 539 567
rect 352 564 539 565
rect 51 559 83 560
rect 51 557 55 559
rect 57 557 80 559
rect 82 557 83 559
rect 51 555 83 557
rect 155 559 187 560
rect 155 557 159 559
rect 161 557 184 559
rect 186 557 187 559
rect 155 555 187 557
rect 302 558 306 559
rect 302 556 303 558
rect 305 556 306 558
rect 7 550 92 551
rect 7 548 89 550
rect 91 548 92 550
rect 7 547 92 548
rect 103 550 219 551
rect 103 548 104 550
rect 106 548 216 550
rect 218 548 219 550
rect 103 547 219 548
rect 7 514 11 547
rect 80 542 115 543
rect 80 540 81 542
rect 83 540 112 542
rect 114 540 115 542
rect 80 539 115 540
rect 206 537 219 538
rect 62 535 75 536
rect 16 533 23 535
rect 16 531 19 533
rect 21 531 23 533
rect 62 533 63 535
rect 65 533 72 535
rect 74 533 75 535
rect 62 532 75 533
rect 166 535 179 536
rect 166 533 167 535
rect 169 533 176 535
rect 178 533 179 535
rect 206 535 208 537
rect 210 535 216 537
rect 218 535 219 537
rect 206 533 219 535
rect 247 533 260 534
rect 166 532 179 533
rect 16 530 23 531
rect 171 527 175 532
rect 247 531 257 533
rect 259 531 260 533
rect 247 530 260 531
rect 247 527 251 530
rect 171 523 251 527
rect 3 510 11 514
rect 7 472 11 510
rect 251 505 255 507
rect 251 503 252 505
rect 254 503 255 505
rect 251 501 255 503
rect 83 491 255 495
rect 83 486 87 491
rect 251 488 255 491
rect 242 486 246 487
rect 79 485 92 486
rect 39 483 52 485
rect 39 481 40 483
rect 42 481 48 483
rect 50 481 52 483
rect 79 483 80 485
rect 82 483 89 485
rect 91 483 92 485
rect 79 482 92 483
rect 183 485 196 486
rect 183 483 184 485
rect 186 483 193 485
rect 195 483 196 485
rect 242 484 243 486
rect 245 484 246 486
rect 242 483 246 484
rect 251 486 260 488
rect 251 484 257 486
rect 259 484 260 486
rect 251 483 260 484
rect 183 482 196 483
rect 39 480 52 481
rect 143 478 178 479
rect 143 476 144 478
rect 146 476 175 478
rect 177 476 178 478
rect 143 475 178 476
rect 7 470 8 472
rect 10 470 11 472
rect 7 469 11 470
rect 39 470 155 471
rect 39 468 40 470
rect 42 468 152 470
rect 154 468 155 470
rect 39 467 155 468
rect 176 470 251 471
rect 176 468 177 470
rect 179 468 251 470
rect 176 467 251 468
rect 71 461 103 463
rect 71 459 72 461
rect 74 459 97 461
rect 99 459 103 461
rect 71 458 103 459
rect 175 461 207 463
rect 175 459 176 461
rect 178 459 201 461
rect 203 459 207 461
rect 175 458 207 459
rect 3 444 7 445
rect 3 442 4 444
rect 6 442 7 444
rect 3 441 7 442
rect 3 434 7 435
rect 3 432 4 434
rect 6 432 7 434
rect 3 431 7 432
rect 51 415 83 416
rect 51 413 55 415
rect 57 413 80 415
rect 82 413 83 415
rect 51 411 83 413
rect 155 415 187 416
rect 155 413 159 415
rect 161 413 184 415
rect 186 413 187 415
rect 155 411 187 413
rect 247 409 251 467
rect 247 407 248 409
rect 250 407 251 409
rect 3 406 92 407
rect 3 404 81 406
rect 83 404 92 406
rect 3 403 92 404
rect 103 406 219 407
rect 103 404 104 406
rect 106 404 216 406
rect 218 404 219 406
rect 247 405 251 407
rect 302 462 306 556
rect 326 558 416 560
rect 326 556 329 558
rect 331 556 361 558
rect 363 556 411 558
rect 413 556 416 558
rect 326 555 416 556
rect 456 558 475 559
rect 456 556 457 558
rect 459 556 472 558
rect 474 556 475 558
rect 456 555 475 556
rect 535 558 539 564
rect 535 556 536 558
rect 538 556 539 558
rect 535 555 539 556
rect 584 558 603 559
rect 584 556 585 558
rect 587 556 600 558
rect 602 556 603 558
rect 584 555 603 556
rect 392 543 500 544
rect 392 541 393 543
rect 395 541 497 543
rect 499 541 500 543
rect 392 540 500 541
rect 560 543 564 544
rect 560 541 561 543
rect 563 541 564 543
rect 560 540 564 541
rect 624 541 628 542
rect 624 539 625 541
rect 627 539 628 541
rect 624 535 628 539
rect 311 534 405 535
rect 311 532 313 534
rect 315 532 321 534
rect 323 533 405 534
rect 323 532 361 533
rect 311 531 361 532
rect 363 531 402 533
rect 404 531 405 533
rect 520 534 628 535
rect 520 532 521 534
rect 523 532 628 534
rect 520 531 628 532
rect 311 530 405 531
rect 464 525 533 526
rect 464 523 466 525
rect 468 523 530 525
rect 532 523 533 525
rect 464 522 533 523
rect 592 525 597 526
rect 592 523 594 525
rect 596 523 597 525
rect 592 522 597 523
rect 464 495 533 496
rect 464 493 465 495
rect 467 493 530 495
rect 532 493 533 495
rect 464 492 533 493
rect 593 495 597 496
rect 593 493 594 495
rect 596 493 597 495
rect 593 492 597 493
rect 311 487 405 488
rect 311 485 313 487
rect 315 485 321 487
rect 323 485 361 487
rect 363 485 402 487
rect 404 485 405 487
rect 311 484 405 485
rect 520 486 628 487
rect 520 484 521 486
rect 523 484 628 486
rect 520 483 628 484
rect 624 479 628 483
rect 392 477 500 478
rect 392 475 393 477
rect 395 475 497 477
rect 499 475 500 477
rect 392 474 500 475
rect 560 477 564 478
rect 560 475 561 477
rect 563 475 564 477
rect 624 477 625 479
rect 627 477 628 479
rect 624 476 628 477
rect 560 474 564 475
rect 302 460 303 462
rect 305 460 306 462
rect 302 414 306 460
rect 327 461 416 463
rect 327 459 329 461
rect 331 459 361 461
rect 363 459 411 461
rect 413 459 416 461
rect 456 462 475 463
rect 456 460 457 462
rect 459 460 472 462
rect 474 460 475 462
rect 456 459 475 460
rect 535 462 539 463
rect 535 460 536 462
rect 538 460 539 462
rect 327 458 416 459
rect 535 454 539 460
rect 584 462 603 463
rect 584 460 585 462
rect 587 460 600 462
rect 602 460 603 462
rect 584 459 603 460
rect 352 453 539 454
rect 352 451 353 453
rect 355 451 539 453
rect 352 450 539 451
rect 352 423 539 424
rect 352 421 353 423
rect 355 421 539 423
rect 352 420 539 421
rect 302 412 303 414
rect 305 412 306 414
rect 103 403 219 404
rect 3 327 7 403
rect 80 398 115 399
rect 80 396 81 398
rect 83 396 112 398
rect 114 396 115 398
rect 80 395 115 396
rect 206 393 219 394
rect 62 391 75 392
rect 17 389 23 390
rect 17 387 19 389
rect 21 387 23 389
rect 62 389 63 391
rect 65 389 72 391
rect 74 389 75 391
rect 62 388 75 389
rect 166 391 179 392
rect 166 389 167 391
rect 169 389 176 391
rect 178 389 179 391
rect 206 391 208 393
rect 210 391 216 393
rect 218 391 219 393
rect 206 389 219 391
rect 251 389 260 390
rect 166 388 179 389
rect 17 386 23 387
rect 171 384 175 388
rect 251 387 257 389
rect 259 387 260 389
rect 251 386 260 387
rect 251 384 255 386
rect 171 380 255 384
rect 251 370 255 373
rect 251 368 252 370
rect 254 368 255 370
rect 251 367 255 368
rect 251 361 255 363
rect 251 359 252 361
rect 254 359 255 361
rect 251 357 255 359
rect 83 348 251 352
rect 83 342 87 348
rect 246 344 251 348
rect 235 343 242 344
rect 79 341 92 342
rect 39 339 52 341
rect 39 337 40 339
rect 42 337 48 339
rect 50 337 52 339
rect 79 339 80 341
rect 82 339 89 341
rect 91 339 92 341
rect 79 338 92 339
rect 183 341 196 342
rect 183 339 184 341
rect 186 339 193 341
rect 195 339 196 341
rect 235 341 237 343
rect 239 341 242 343
rect 235 339 242 341
rect 246 342 260 344
rect 246 340 257 342
rect 259 340 260 342
rect 246 339 260 340
rect 183 338 196 339
rect 39 336 52 337
rect 143 334 178 335
rect 143 332 144 334
rect 146 332 175 334
rect 177 332 178 334
rect 143 331 178 332
rect 3 326 11 327
rect 3 324 8 326
rect 10 324 11 326
rect 3 323 11 324
rect 39 326 155 327
rect 39 324 40 326
rect 42 324 152 326
rect 154 324 155 326
rect 39 323 155 324
rect 302 319 306 412
rect 327 414 416 416
rect 327 412 329 414
rect 331 412 361 414
rect 363 412 412 414
rect 414 412 416 414
rect 327 411 416 412
rect 456 414 475 415
rect 456 412 457 414
rect 459 412 472 414
rect 474 412 475 414
rect 456 411 475 412
rect 535 414 539 420
rect 535 412 536 414
rect 538 412 539 414
rect 535 411 539 412
rect 584 414 603 415
rect 584 412 585 414
rect 587 412 600 414
rect 602 412 603 414
rect 584 411 603 412
rect 392 399 500 400
rect 392 397 393 399
rect 395 397 497 399
rect 499 397 500 399
rect 392 396 500 397
rect 560 398 564 399
rect 560 396 561 398
rect 563 396 564 398
rect 560 395 564 396
rect 624 397 628 398
rect 624 395 625 397
rect 627 395 628 397
rect 624 391 628 395
rect 311 389 405 391
rect 311 387 312 389
rect 314 387 321 389
rect 323 387 361 389
rect 363 387 401 389
rect 403 387 405 389
rect 520 390 628 391
rect 520 388 521 390
rect 523 388 628 390
rect 520 387 628 388
rect 311 386 405 387
rect 464 381 533 382
rect 464 379 465 381
rect 467 379 530 381
rect 532 379 533 381
rect 464 378 533 379
rect 593 381 597 382
rect 593 379 594 381
rect 596 379 597 381
rect 593 378 597 379
rect 464 351 533 352
rect 464 349 465 351
rect 467 349 530 351
rect 532 349 533 351
rect 464 348 533 349
rect 593 351 597 352
rect 593 349 594 351
rect 596 349 597 351
rect 593 348 597 349
rect 311 342 405 344
rect 311 340 312 342
rect 314 340 321 342
rect 323 340 361 342
rect 363 340 401 342
rect 403 340 405 342
rect 311 338 405 340
rect 520 342 628 343
rect 520 340 521 342
rect 523 340 628 342
rect 520 339 628 340
rect 624 335 628 339
rect 392 333 500 334
rect 392 331 393 333
rect 395 331 497 333
rect 499 331 500 333
rect 392 330 500 331
rect 560 333 564 334
rect 560 331 561 333
rect 563 331 564 333
rect 624 333 625 335
rect 627 333 628 335
rect 624 332 628 333
rect 560 330 564 331
rect 71 317 103 319
rect 71 315 72 317
rect 74 315 97 317
rect 99 315 103 317
rect 71 314 103 315
rect 175 317 251 319
rect 175 315 176 317
rect 178 315 201 317
rect 203 315 251 317
rect 175 314 251 315
rect 295 317 306 319
rect 295 315 303 317
rect 305 315 306 317
rect 295 314 306 315
rect 327 318 416 319
rect 327 316 329 318
rect 331 317 413 318
rect 331 316 361 317
rect 327 315 361 316
rect 363 316 413 317
rect 415 316 416 318
rect 363 315 416 316
rect 456 318 475 319
rect 456 316 457 318
rect 459 316 472 318
rect 474 316 475 318
rect 456 315 475 316
rect 535 318 539 319
rect 535 316 536 318
rect 538 316 539 318
rect 327 314 416 315
rect 3 298 7 299
rect 3 296 4 298
rect 6 296 7 298
rect 3 295 7 296
rect 3 290 7 291
rect 3 288 4 290
rect 6 288 7 290
rect 3 287 7 288
rect 51 271 83 272
rect 51 269 55 271
rect 57 269 80 271
rect 82 269 83 271
rect 51 267 83 269
rect 155 271 187 272
rect 155 269 159 271
rect 161 269 184 271
rect 186 269 187 271
rect 155 267 187 269
rect 7 262 92 263
rect 7 260 89 262
rect 91 260 92 262
rect 7 259 92 260
rect 103 262 219 263
rect 103 260 104 262
rect 106 260 216 262
rect 218 260 219 262
rect 103 259 219 260
rect 247 259 251 314
rect 7 226 11 259
rect 247 257 248 259
rect 250 257 251 259
rect 247 255 251 257
rect 302 270 306 314
rect 535 310 539 316
rect 584 318 603 319
rect 584 316 585 318
rect 587 316 600 318
rect 602 316 603 318
rect 584 315 603 316
rect 352 309 539 310
rect 352 307 353 309
rect 355 307 539 309
rect 352 306 539 307
rect 352 279 539 280
rect 352 277 353 279
rect 355 277 539 279
rect 352 276 539 277
rect 302 268 303 270
rect 305 268 306 270
rect 80 254 115 255
rect 80 252 81 254
rect 83 252 112 254
rect 114 252 115 254
rect 80 251 115 252
rect 206 249 219 250
rect 62 247 75 248
rect 16 245 23 247
rect 16 243 19 245
rect 21 243 23 245
rect 62 245 63 247
rect 65 245 72 247
rect 74 245 75 247
rect 62 244 75 245
rect 166 247 179 248
rect 166 245 167 247
rect 169 245 176 247
rect 178 245 179 247
rect 206 247 208 249
rect 210 247 216 249
rect 218 247 219 249
rect 206 245 219 247
rect 247 245 260 246
rect 166 244 179 245
rect 16 242 23 243
rect 171 239 175 244
rect 247 243 257 245
rect 259 243 260 245
rect 247 242 260 243
rect 247 239 251 242
rect 171 235 251 239
rect 3 222 11 226
rect 251 227 255 229
rect 251 225 252 227
rect 254 225 255 227
rect 251 223 255 225
rect 7 184 11 222
rect 251 217 255 219
rect 251 215 252 217
rect 254 215 255 217
rect 251 213 255 215
rect 83 203 255 207
rect 83 198 87 203
rect 251 200 255 203
rect 242 198 246 199
rect 79 197 92 198
rect 39 195 52 197
rect 39 193 40 195
rect 42 193 48 195
rect 50 193 52 195
rect 79 195 80 197
rect 82 195 89 197
rect 91 195 92 197
rect 79 194 92 195
rect 183 197 196 198
rect 183 195 184 197
rect 186 195 193 197
rect 195 195 196 197
rect 242 196 243 198
rect 245 196 246 198
rect 242 195 246 196
rect 251 198 260 200
rect 251 196 257 198
rect 259 196 260 198
rect 251 195 260 196
rect 183 194 196 195
rect 39 192 52 193
rect 143 190 178 191
rect 143 188 144 190
rect 146 188 175 190
rect 177 188 178 190
rect 143 187 178 188
rect 7 182 8 184
rect 10 182 11 184
rect 7 181 11 182
rect 39 182 155 183
rect 39 180 40 182
rect 42 180 152 182
rect 154 180 155 182
rect 39 179 155 180
rect 176 182 251 183
rect 176 180 177 182
rect 179 180 251 182
rect 176 179 251 180
rect 71 173 103 175
rect 71 171 72 173
rect 74 171 97 173
rect 99 171 103 173
rect 71 170 103 171
rect 175 173 207 175
rect 175 171 176 173
rect 178 171 201 173
rect 203 171 207 173
rect 175 170 207 171
rect 3 156 7 157
rect 3 154 4 156
rect 6 154 7 156
rect 3 153 7 154
rect 3 146 7 147
rect 3 144 4 146
rect 6 144 7 146
rect 3 143 7 144
rect 51 127 83 128
rect 51 125 55 127
rect 57 125 80 127
rect 82 125 83 127
rect 51 123 83 125
rect 155 127 187 128
rect 155 125 159 127
rect 161 125 184 127
rect 186 125 187 127
rect 155 123 187 125
rect 247 120 251 179
rect 3 118 92 119
rect 3 116 81 118
rect 83 116 92 118
rect 3 115 92 116
rect 103 118 219 119
rect 103 116 104 118
rect 106 116 216 118
rect 218 116 219 118
rect 247 118 248 120
rect 250 118 251 120
rect 247 117 251 118
rect 302 174 306 268
rect 326 271 416 272
rect 326 269 329 271
rect 331 270 412 271
rect 331 269 361 270
rect 326 268 361 269
rect 363 269 412 270
rect 414 269 416 271
rect 363 268 416 269
rect 326 267 416 268
rect 456 270 475 271
rect 456 268 457 270
rect 459 268 472 270
rect 474 268 475 270
rect 456 267 475 268
rect 535 270 539 276
rect 535 268 536 270
rect 538 268 539 270
rect 535 267 539 268
rect 584 270 603 271
rect 584 268 585 270
rect 587 268 600 270
rect 602 268 603 270
rect 584 267 603 268
rect 392 255 500 256
rect 392 253 393 255
rect 395 253 497 255
rect 499 253 500 255
rect 392 252 500 253
rect 560 255 564 256
rect 560 253 561 255
rect 563 253 564 255
rect 560 252 564 253
rect 624 253 628 254
rect 624 251 625 253
rect 627 251 628 253
rect 624 247 628 251
rect 311 245 405 247
rect 311 243 312 245
rect 314 243 321 245
rect 323 243 361 245
rect 363 243 401 245
rect 403 243 405 245
rect 520 246 628 247
rect 520 244 521 246
rect 523 244 628 246
rect 520 243 628 244
rect 311 242 405 243
rect 464 237 533 238
rect 464 235 465 237
rect 467 235 529 237
rect 531 235 533 237
rect 464 234 533 235
rect 593 237 597 238
rect 593 235 594 237
rect 596 235 597 237
rect 593 234 597 235
rect 464 207 533 208
rect 464 205 465 207
rect 467 205 529 207
rect 531 205 533 207
rect 464 204 533 205
rect 593 207 597 208
rect 593 205 594 207
rect 596 205 597 207
rect 593 204 597 205
rect 311 198 405 200
rect 311 196 312 198
rect 314 196 321 198
rect 323 196 361 198
rect 363 196 401 198
rect 403 196 405 198
rect 311 195 405 196
rect 520 198 628 199
rect 520 196 521 198
rect 523 196 628 198
rect 520 195 628 196
rect 624 191 628 195
rect 392 189 500 190
rect 392 187 393 189
rect 395 187 497 189
rect 499 187 500 189
rect 392 186 500 187
rect 560 189 564 190
rect 560 187 561 189
rect 563 187 564 189
rect 624 189 625 191
rect 627 189 628 191
rect 624 188 628 189
rect 560 186 564 187
rect 302 172 303 174
rect 305 172 306 174
rect 302 126 306 172
rect 327 174 416 175
rect 327 173 412 174
rect 327 171 329 173
rect 331 171 361 173
rect 363 172 412 173
rect 414 172 416 174
rect 363 171 416 172
rect 456 174 475 175
rect 456 172 457 174
rect 459 172 472 174
rect 474 172 475 174
rect 456 171 475 172
rect 535 174 539 175
rect 535 172 536 174
rect 538 172 539 174
rect 327 170 416 171
rect 535 166 539 172
rect 584 174 603 175
rect 584 172 585 174
rect 587 172 600 174
rect 602 172 603 174
rect 584 171 603 172
rect 352 165 539 166
rect 352 163 353 165
rect 355 163 539 165
rect 352 162 539 163
rect 352 135 539 136
rect 352 133 353 135
rect 355 133 539 135
rect 352 132 539 133
rect 302 124 303 126
rect 305 124 306 126
rect 103 115 219 116
rect 3 39 7 115
rect 80 110 115 111
rect 80 108 81 110
rect 83 108 112 110
rect 114 108 115 110
rect 80 107 115 108
rect 206 105 219 106
rect 62 103 75 104
rect 18 101 23 103
rect 18 99 19 101
rect 21 99 23 101
rect 62 101 63 103
rect 65 101 72 103
rect 74 101 75 103
rect 62 100 75 101
rect 166 103 179 104
rect 166 101 167 103
rect 169 101 176 103
rect 178 101 179 103
rect 206 103 208 105
rect 210 103 216 105
rect 218 103 219 105
rect 206 101 219 103
rect 251 101 260 102
rect 166 100 179 101
rect 18 98 23 99
rect 171 96 175 100
rect 251 99 257 101
rect 259 99 260 101
rect 251 98 260 99
rect 251 96 255 98
rect 171 92 255 96
rect 251 82 255 85
rect 251 80 252 82
rect 254 80 255 82
rect 251 79 255 80
rect 83 60 251 64
rect 83 54 87 60
rect 246 56 251 60
rect 246 54 260 56
rect 79 53 92 54
rect 39 51 52 53
rect 39 49 40 51
rect 42 49 48 51
rect 50 49 52 51
rect 79 51 80 53
rect 82 51 89 53
rect 91 51 92 53
rect 79 50 92 51
rect 183 53 196 54
rect 183 51 184 53
rect 186 51 193 53
rect 195 51 196 53
rect 246 52 257 54
rect 259 52 260 54
rect 246 51 260 52
rect 183 50 196 51
rect 39 48 52 49
rect 143 46 178 47
rect 143 44 144 46
rect 146 44 175 46
rect 177 44 178 46
rect 143 43 178 44
rect 247 45 251 46
rect 247 43 248 45
rect 250 43 251 45
rect 247 42 251 43
rect 3 38 11 39
rect 3 36 8 38
rect 10 36 11 38
rect 3 35 11 36
rect 39 38 155 39
rect 39 36 40 38
rect 42 36 152 38
rect 154 36 155 38
rect 39 35 155 36
rect 302 31 306 124
rect 327 127 416 128
rect 327 126 361 127
rect 327 124 329 126
rect 331 125 361 126
rect 363 125 412 127
rect 414 125 416 127
rect 331 124 416 125
rect 327 123 416 124
rect 456 126 475 127
rect 456 124 457 126
rect 459 124 472 126
rect 474 124 475 126
rect 456 123 475 124
rect 535 126 539 132
rect 535 124 536 126
rect 538 124 539 126
rect 535 123 539 124
rect 584 126 603 127
rect 584 124 585 126
rect 587 124 600 126
rect 602 124 603 126
rect 584 123 603 124
rect 392 110 500 111
rect 392 108 393 110
rect 395 108 497 110
rect 499 108 500 110
rect 392 107 500 108
rect 560 110 564 111
rect 560 108 561 110
rect 563 108 564 110
rect 560 107 564 108
rect 624 109 628 110
rect 624 107 625 109
rect 627 107 628 109
rect 624 103 628 107
rect 311 101 405 103
rect 311 99 312 101
rect 314 99 321 101
rect 323 99 361 101
rect 363 99 401 101
rect 403 99 405 101
rect 520 102 628 103
rect 520 100 521 102
rect 523 100 628 102
rect 520 99 628 100
rect 311 98 405 99
rect 464 93 533 94
rect 464 91 465 93
rect 467 91 529 93
rect 531 91 533 93
rect 464 90 533 91
rect 593 93 597 94
rect 593 91 594 93
rect 596 91 597 93
rect 593 90 597 91
rect 464 63 533 64
rect 464 61 465 63
rect 467 61 530 63
rect 532 61 533 63
rect 464 60 533 61
rect 592 63 597 64
rect 592 61 594 63
rect 596 61 597 63
rect 592 60 597 61
rect 311 55 405 56
rect 311 54 361 55
rect 311 52 312 54
rect 314 52 321 54
rect 323 53 361 54
rect 363 54 405 55
rect 363 53 401 54
rect 323 52 401 53
rect 403 52 405 54
rect 311 51 405 52
rect 520 54 628 55
rect 520 52 521 54
rect 523 52 628 54
rect 520 51 628 52
rect 624 47 628 51
rect 392 45 500 46
rect 392 43 393 45
rect 395 43 497 45
rect 499 43 500 45
rect 392 42 500 43
rect 560 45 564 46
rect 560 43 561 45
rect 563 43 564 45
rect 624 45 625 47
rect 627 45 628 47
rect 624 44 628 45
rect 560 42 564 43
rect 71 29 103 31
rect 71 27 72 29
rect 74 27 97 29
rect 99 27 103 29
rect 71 26 103 27
rect 175 29 306 31
rect 175 27 176 29
rect 178 27 201 29
rect 203 27 303 29
rect 305 27 306 29
rect 175 26 306 27
rect 327 30 416 31
rect 327 29 412 30
rect 327 27 329 29
rect 331 27 361 29
rect 363 28 412 29
rect 414 28 416 30
rect 363 27 416 28
rect 456 30 484 31
rect 456 28 457 30
rect 459 28 478 30
rect 480 28 484 30
rect 456 27 484 28
rect 535 30 539 31
rect 535 28 536 30
rect 538 28 539 30
rect 327 26 416 27
rect 96 22 101 26
rect 327 22 332 26
rect 535 22 539 28
rect 584 30 603 31
rect 584 28 585 30
rect 587 28 600 30
rect 602 28 603 30
rect 584 27 603 28
rect 96 17 332 22
rect 352 21 539 22
rect 352 19 353 21
rect 355 19 539 21
rect 352 18 539 19
rect 3 10 7 11
rect 3 8 4 10
rect 6 8 7 10
rect 3 7 7 8
<< alu3 >>
rect 3 578 7 579
rect 3 576 4 578
rect 6 576 7 578
rect 3 444 7 576
rect 182 559 187 560
rect 182 557 184 559
rect 186 557 187 559
rect 182 555 187 557
rect 327 558 332 560
rect 327 556 329 558
rect 331 556 332 558
rect 327 555 332 556
rect 560 543 564 544
rect 560 541 561 543
rect 563 541 564 543
rect 560 540 564 541
rect 16 533 23 535
rect 16 531 19 533
rect 21 531 23 533
rect 16 530 23 531
rect 464 525 469 526
rect 464 523 466 525
rect 468 523 469 525
rect 464 522 469 523
rect 592 525 597 526
rect 592 523 594 525
rect 596 523 597 525
rect 592 522 597 523
rect 251 505 255 507
rect 251 503 252 505
rect 254 503 255 505
rect 242 486 246 487
rect 242 484 243 486
rect 245 484 246 486
rect 242 483 246 484
rect 95 461 103 463
rect 95 459 97 461
rect 99 459 103 461
rect 95 458 103 459
rect 3 442 4 444
rect 6 442 7 444
rect 3 441 7 442
rect 3 434 7 435
rect 3 432 4 434
rect 6 432 7 434
rect 3 298 7 432
rect 182 415 187 416
rect 182 413 184 415
rect 186 413 187 415
rect 182 411 187 413
rect 17 389 23 390
rect 17 387 19 389
rect 21 387 23 389
rect 17 386 23 387
rect 251 370 255 503
rect 464 495 468 522
rect 464 493 465 495
rect 467 493 468 495
rect 327 461 332 463
rect 327 459 329 461
rect 331 459 332 461
rect 327 458 332 459
rect 327 414 332 416
rect 327 412 329 414
rect 331 412 332 414
rect 327 411 332 412
rect 251 368 252 370
rect 254 368 255 370
rect 251 367 255 368
rect 464 381 468 493
rect 593 495 597 522
rect 593 493 594 495
rect 596 493 597 495
rect 560 477 564 478
rect 560 475 561 477
rect 563 475 564 477
rect 560 474 564 475
rect 560 398 564 399
rect 560 396 561 398
rect 563 396 564 398
rect 560 395 564 396
rect 464 379 465 381
rect 467 379 468 381
rect 251 361 255 363
rect 251 359 252 361
rect 254 359 255 361
rect 235 343 242 344
rect 235 341 237 343
rect 239 341 242 343
rect 235 339 242 341
rect 95 317 103 319
rect 95 315 97 317
rect 99 315 103 317
rect 95 314 103 315
rect 3 296 4 298
rect 6 296 7 298
rect 3 295 7 296
rect 3 290 7 291
rect 3 288 4 290
rect 6 288 7 290
rect 3 156 7 288
rect 155 271 163 272
rect 155 269 159 271
rect 161 269 163 271
rect 155 267 163 269
rect 16 245 23 247
rect 16 243 19 245
rect 21 243 23 245
rect 16 242 23 243
rect 251 227 255 359
rect 464 351 468 379
rect 464 349 465 351
rect 467 349 468 351
rect 327 318 332 319
rect 327 316 329 318
rect 331 316 332 318
rect 327 314 332 316
rect 327 271 332 272
rect 327 269 329 271
rect 331 269 332 271
rect 327 267 332 269
rect 251 225 252 227
rect 254 225 255 227
rect 251 223 255 225
rect 464 238 468 349
rect 593 381 597 493
rect 593 379 594 381
rect 596 379 597 381
rect 593 351 597 379
rect 593 349 594 351
rect 596 349 597 351
rect 560 333 564 334
rect 560 331 561 333
rect 563 331 564 333
rect 560 330 564 331
rect 560 255 564 256
rect 560 253 561 255
rect 563 253 564 255
rect 560 252 564 253
rect 464 237 469 238
rect 464 235 465 237
rect 467 235 469 237
rect 464 234 469 235
rect 593 237 597 349
rect 593 235 594 237
rect 596 235 597 237
rect 251 217 255 219
rect 251 215 252 217
rect 254 215 255 217
rect 242 198 246 199
rect 242 196 243 198
rect 245 196 246 198
rect 242 195 246 196
rect 95 173 103 175
rect 95 171 97 173
rect 99 171 103 173
rect 95 170 103 171
rect 3 154 4 156
rect 6 154 7 156
rect 3 153 7 154
rect 3 146 7 147
rect 3 144 4 146
rect 6 144 7 146
rect 3 10 7 144
rect 158 127 163 128
rect 158 125 159 127
rect 161 125 163 127
rect 158 123 163 125
rect 18 101 23 103
rect 18 99 19 101
rect 21 99 23 101
rect 18 98 23 99
rect 251 82 255 215
rect 464 207 468 234
rect 464 205 465 207
rect 467 205 468 207
rect 327 173 332 175
rect 327 171 329 173
rect 331 171 332 173
rect 327 170 332 171
rect 327 126 332 128
rect 327 124 329 126
rect 331 124 332 126
rect 327 123 332 124
rect 251 80 252 82
rect 254 80 255 82
rect 251 79 255 80
rect 464 94 468 205
rect 593 207 597 235
rect 593 205 594 207
rect 596 205 597 207
rect 560 189 564 190
rect 560 187 561 189
rect 563 187 564 189
rect 560 186 564 187
rect 560 110 564 111
rect 560 108 561 110
rect 563 108 564 110
rect 560 107 564 108
rect 464 93 469 94
rect 464 91 465 93
rect 467 91 469 93
rect 464 90 469 91
rect 593 93 597 205
rect 593 91 594 93
rect 596 91 597 93
rect 464 63 468 90
rect 593 64 597 91
rect 464 61 465 63
rect 467 61 468 63
rect 464 60 468 61
rect 592 63 597 64
rect 592 61 594 63
rect 596 61 597 63
rect 592 60 597 61
rect 247 45 564 46
rect 247 43 248 45
rect 250 43 561 45
rect 563 43 564 45
rect 247 42 564 43
rect 3 8 4 10
rect 6 8 7 10
rect 3 7 7 8
<< alu4 >>
rect 182 559 332 560
rect 182 557 184 559
rect 186 558 332 559
rect 186 557 329 558
rect 182 556 329 557
rect 331 556 332 558
rect 182 555 332 556
rect 16 543 564 544
rect 16 541 561 543
rect 563 541 564 543
rect 16 540 564 541
rect 16 535 20 540
rect 16 533 23 535
rect 16 531 19 533
rect 21 531 23 533
rect 16 530 23 531
rect 242 486 564 487
rect 242 484 243 486
rect 245 484 564 486
rect 242 483 564 484
rect 560 477 564 483
rect 560 475 561 477
rect 563 475 564 477
rect 560 474 564 475
rect 95 461 332 463
rect 95 459 97 461
rect 99 459 329 461
rect 331 459 332 461
rect 95 458 332 459
rect 182 415 332 416
rect 182 413 184 415
rect 186 414 332 415
rect 186 413 329 414
rect 182 412 329 413
rect 331 412 332 414
rect 182 411 332 412
rect 560 398 564 400
rect 560 396 561 398
rect 563 396 564 398
rect 560 390 564 396
rect 17 389 564 390
rect 17 387 19 389
rect 21 387 564 389
rect 17 386 564 387
rect 235 343 564 344
rect 235 341 237 343
rect 239 341 564 343
rect 235 340 564 341
rect 235 339 242 340
rect 560 333 564 340
rect 560 331 561 333
rect 563 331 564 333
rect 560 330 564 331
rect 95 318 332 319
rect 95 317 329 318
rect 95 315 97 317
rect 99 316 329 317
rect 331 316 332 318
rect 99 315 332 316
rect 95 314 332 315
rect 155 271 332 272
rect 155 269 159 271
rect 161 269 329 271
rect 331 269 332 271
rect 155 267 332 269
rect 16 255 564 256
rect 16 253 561 255
rect 563 253 564 255
rect 16 252 564 253
rect 16 247 20 252
rect 560 250 564 252
rect 16 245 23 247
rect 16 243 19 245
rect 21 243 23 245
rect 16 242 23 243
rect 242 198 564 200
rect 242 196 243 198
rect 245 196 564 198
rect 242 195 247 196
rect 560 189 564 196
rect 560 187 561 189
rect 563 187 564 189
rect 560 186 564 187
rect 95 173 332 175
rect 95 171 97 173
rect 99 171 329 173
rect 331 171 332 173
rect 95 170 332 171
rect 158 127 332 128
rect 158 125 159 127
rect 161 126 332 127
rect 161 125 329 126
rect 158 124 329 125
rect 331 124 332 126
rect 158 123 332 124
rect 18 110 564 111
rect 18 108 561 110
rect 563 108 564 110
rect 18 107 564 108
rect 18 101 23 107
rect 18 99 19 101
rect 21 99 23 101
rect 18 98 23 99
<< ptie >>
rect 60 576 66 578
rect 60 574 62 576
rect 64 574 66 576
rect 60 572 66 574
rect 100 576 106 578
rect 100 574 102 576
rect 104 574 106 576
rect 100 572 106 574
rect 164 576 170 578
rect 164 574 166 576
rect 168 574 170 576
rect 164 572 170 574
rect 204 576 210 578
rect 204 574 206 576
rect 208 574 210 576
rect 244 576 250 578
rect 244 574 246 576
rect 248 574 250 576
rect 204 572 210 574
rect 244 572 250 574
rect 309 576 315 578
rect 309 574 311 576
rect 313 574 315 576
rect 309 572 315 574
rect 349 576 355 578
rect 349 574 351 576
rect 353 574 355 576
rect 389 576 395 578
rect 389 574 391 576
rect 393 574 395 576
rect 349 572 355 574
rect 389 572 395 574
rect 401 576 407 578
rect 401 574 403 576
rect 405 574 407 576
rect 401 572 407 574
rect 8 444 14 446
rect 48 444 54 446
rect 8 442 10 444
rect 12 442 14 444
rect 8 440 14 442
rect 48 442 50 444
rect 52 442 54 444
rect 48 440 54 442
rect 88 444 94 446
rect 88 442 90 444
rect 92 442 94 444
rect 88 440 94 442
rect 152 444 158 446
rect 152 442 154 444
rect 156 442 158 444
rect 152 440 158 442
rect 192 444 198 446
rect 192 442 194 444
rect 196 442 198 444
rect 192 440 198 442
rect 309 444 315 446
rect 309 442 311 444
rect 313 442 315 444
rect 309 440 315 442
rect 349 444 355 446
rect 389 444 395 446
rect 349 442 351 444
rect 353 442 355 444
rect 349 440 355 442
rect 389 442 391 444
rect 393 442 395 444
rect 389 440 395 442
rect 401 444 407 446
rect 401 442 403 444
rect 405 442 407 444
rect 401 440 407 442
rect 60 432 66 434
rect 60 430 62 432
rect 64 430 66 432
rect 60 428 66 430
rect 100 432 106 434
rect 100 430 102 432
rect 104 430 106 432
rect 100 428 106 430
rect 164 432 170 434
rect 164 430 166 432
rect 168 430 170 432
rect 164 428 170 430
rect 204 432 210 434
rect 204 430 206 432
rect 208 430 210 432
rect 244 432 250 434
rect 244 430 246 432
rect 248 430 250 432
rect 204 428 210 430
rect 244 428 250 430
rect 309 432 315 434
rect 309 430 311 432
rect 313 430 315 432
rect 309 428 315 430
rect 349 432 355 434
rect 349 430 351 432
rect 353 430 355 432
rect 389 432 395 434
rect 389 430 391 432
rect 393 430 395 432
rect 349 428 355 430
rect 389 428 395 430
rect 401 432 407 434
rect 401 430 403 432
rect 405 430 407 432
rect 401 428 407 430
rect 8 300 14 302
rect 48 300 54 302
rect 8 298 10 300
rect 12 298 14 300
rect 8 296 14 298
rect 48 298 50 300
rect 52 298 54 300
rect 48 296 54 298
rect 88 300 94 302
rect 88 298 90 300
rect 92 298 94 300
rect 88 296 94 298
rect 152 300 158 302
rect 152 298 154 300
rect 156 298 158 300
rect 152 296 158 298
rect 192 300 198 302
rect 192 298 194 300
rect 196 298 198 300
rect 192 296 198 298
rect 309 300 315 302
rect 309 298 311 300
rect 313 298 315 300
rect 309 296 315 298
rect 349 300 355 302
rect 389 300 395 302
rect 349 298 351 300
rect 353 298 355 300
rect 349 296 355 298
rect 389 298 391 300
rect 393 298 395 300
rect 389 296 395 298
rect 401 300 407 302
rect 401 298 403 300
rect 405 298 407 300
rect 401 296 407 298
rect 60 288 66 290
rect 60 286 62 288
rect 64 286 66 288
rect 60 284 66 286
rect 100 288 106 290
rect 100 286 102 288
rect 104 286 106 288
rect 100 284 106 286
rect 164 288 170 290
rect 164 286 166 288
rect 168 286 170 288
rect 164 284 170 286
rect 204 288 210 290
rect 204 286 206 288
rect 208 286 210 288
rect 244 288 250 290
rect 244 286 246 288
rect 248 286 250 288
rect 204 284 210 286
rect 244 284 250 286
rect 309 288 315 290
rect 309 286 311 288
rect 313 286 315 288
rect 309 284 315 286
rect 349 288 355 290
rect 349 286 351 288
rect 353 286 355 288
rect 389 288 395 290
rect 389 286 391 288
rect 393 286 395 288
rect 349 284 355 286
rect 389 284 395 286
rect 401 288 407 290
rect 401 286 403 288
rect 405 286 407 288
rect 401 284 407 286
rect 8 156 14 158
rect 48 156 54 158
rect 8 154 10 156
rect 12 154 14 156
rect 8 152 14 154
rect 48 154 50 156
rect 52 154 54 156
rect 48 152 54 154
rect 88 156 94 158
rect 88 154 90 156
rect 92 154 94 156
rect 88 152 94 154
rect 152 156 158 158
rect 152 154 154 156
rect 156 154 158 156
rect 152 152 158 154
rect 192 156 198 158
rect 192 154 194 156
rect 196 154 198 156
rect 192 152 198 154
rect 309 156 315 158
rect 309 154 311 156
rect 313 154 315 156
rect 309 152 315 154
rect 349 156 355 158
rect 389 156 395 158
rect 349 154 351 156
rect 353 154 355 156
rect 349 152 355 154
rect 389 154 391 156
rect 393 154 395 156
rect 389 152 395 154
rect 401 156 407 158
rect 401 154 403 156
rect 405 154 407 156
rect 401 152 407 154
rect 60 144 66 146
rect 60 142 62 144
rect 64 142 66 144
rect 60 140 66 142
rect 100 144 106 146
rect 100 142 102 144
rect 104 142 106 144
rect 100 140 106 142
rect 164 144 170 146
rect 164 142 166 144
rect 168 142 170 144
rect 164 140 170 142
rect 204 144 210 146
rect 204 142 206 144
rect 208 142 210 144
rect 244 144 250 146
rect 244 142 246 144
rect 248 142 250 144
rect 204 140 210 142
rect 244 140 250 142
rect 309 144 315 146
rect 309 142 311 144
rect 313 142 315 144
rect 309 140 315 142
rect 349 144 355 146
rect 349 142 351 144
rect 353 142 355 144
rect 389 144 395 146
rect 389 142 391 144
rect 393 142 395 144
rect 349 140 355 142
rect 389 140 395 142
rect 401 144 407 146
rect 401 142 403 144
rect 405 142 407 144
rect 401 140 407 142
rect 8 12 14 14
rect 48 12 54 14
rect 8 10 10 12
rect 12 10 14 12
rect 8 8 14 10
rect 48 10 50 12
rect 52 10 54 12
rect 48 8 54 10
rect 88 12 94 14
rect 88 10 90 12
rect 92 10 94 12
rect 88 8 94 10
rect 152 12 158 14
rect 152 10 154 12
rect 156 10 158 12
rect 152 8 158 10
rect 192 12 198 14
rect 192 10 194 12
rect 196 10 198 12
rect 192 8 198 10
rect 309 12 315 14
rect 309 10 311 12
rect 313 10 315 12
rect 309 8 315 10
rect 349 12 355 14
rect 389 12 395 14
rect 349 10 351 12
rect 353 10 355 12
rect 349 8 355 10
rect 389 10 391 12
rect 393 10 395 12
rect 389 8 395 10
rect 401 12 407 14
rect 401 10 403 12
rect 405 10 407 12
rect 401 8 407 10
<< ntie >>
rect 27 516 33 518
rect 27 514 29 516
rect 31 514 33 516
rect 100 516 106 518
rect 27 512 33 514
rect 100 514 102 516
rect 104 514 106 516
rect 131 516 137 518
rect 100 512 106 514
rect 131 514 133 516
rect 135 514 137 516
rect 204 516 210 518
rect 131 512 137 514
rect 204 514 206 516
rect 208 514 210 516
rect 244 516 250 518
rect 204 512 210 514
rect 244 514 246 516
rect 248 514 250 516
rect 276 516 282 518
rect 244 512 250 514
rect 276 514 278 516
rect 280 514 282 516
rect 349 516 355 518
rect 276 512 282 514
rect 349 514 351 516
rect 353 514 355 516
rect 389 516 395 518
rect 349 512 355 514
rect 389 514 391 516
rect 393 514 395 516
rect 434 516 440 518
rect 389 512 395 514
rect 434 514 436 516
rect 438 514 440 516
rect 434 512 440 514
rect 8 504 14 506
rect 8 502 10 504
rect 12 502 14 504
rect 48 504 54 506
rect 8 500 14 502
rect 48 502 50 504
rect 52 502 54 504
rect 121 504 127 506
rect 48 500 54 502
rect 121 502 123 504
rect 125 502 127 504
rect 152 504 158 506
rect 121 500 127 502
rect 152 502 154 504
rect 156 502 158 504
rect 225 504 231 506
rect 152 500 158 502
rect 225 502 227 504
rect 229 502 231 504
rect 276 504 282 506
rect 225 500 231 502
rect 276 502 278 504
rect 280 502 282 504
rect 349 504 355 506
rect 276 500 282 502
rect 349 502 351 504
rect 353 502 355 504
rect 389 504 395 506
rect 349 500 355 502
rect 389 502 391 504
rect 393 502 395 504
rect 434 504 440 506
rect 389 500 395 502
rect 434 502 436 504
rect 438 502 440 504
rect 434 500 440 502
rect 27 372 33 374
rect 27 370 29 372
rect 31 370 33 372
rect 100 372 106 374
rect 27 368 33 370
rect 100 370 102 372
rect 104 370 106 372
rect 131 372 137 374
rect 100 368 106 370
rect 131 370 133 372
rect 135 370 137 372
rect 204 372 210 374
rect 131 368 137 370
rect 204 370 206 372
rect 208 370 210 372
rect 244 372 250 374
rect 204 368 210 370
rect 244 370 246 372
rect 248 370 250 372
rect 276 372 282 374
rect 244 368 250 370
rect 276 370 278 372
rect 280 370 282 372
rect 349 372 355 374
rect 276 368 282 370
rect 349 370 351 372
rect 353 370 355 372
rect 389 372 395 374
rect 349 368 355 370
rect 389 370 391 372
rect 393 370 395 372
rect 434 372 440 374
rect 389 368 395 370
rect 434 370 436 372
rect 438 370 440 372
rect 434 368 440 370
rect 8 360 14 362
rect 8 358 10 360
rect 12 358 14 360
rect 48 360 54 362
rect 8 356 14 358
rect 48 358 50 360
rect 52 358 54 360
rect 121 360 127 362
rect 48 356 54 358
rect 121 358 123 360
rect 125 358 127 360
rect 152 360 158 362
rect 121 356 127 358
rect 152 358 154 360
rect 156 358 158 360
rect 225 360 231 362
rect 152 356 158 358
rect 225 358 227 360
rect 229 358 231 360
rect 276 360 282 362
rect 225 356 231 358
rect 276 358 278 360
rect 280 358 282 360
rect 349 360 355 362
rect 276 356 282 358
rect 349 358 351 360
rect 353 358 355 360
rect 389 360 395 362
rect 349 356 355 358
rect 389 358 391 360
rect 393 358 395 360
rect 434 360 440 362
rect 389 356 395 358
rect 434 358 436 360
rect 438 358 440 360
rect 434 356 440 358
rect 27 228 33 230
rect 27 226 29 228
rect 31 226 33 228
rect 100 228 106 230
rect 27 224 33 226
rect 100 226 102 228
rect 104 226 106 228
rect 131 228 137 230
rect 100 224 106 226
rect 131 226 133 228
rect 135 226 137 228
rect 204 228 210 230
rect 131 224 137 226
rect 204 226 206 228
rect 208 226 210 228
rect 244 228 250 230
rect 204 224 210 226
rect 244 226 246 228
rect 248 226 250 228
rect 276 228 282 230
rect 244 224 250 226
rect 276 226 278 228
rect 280 226 282 228
rect 349 228 355 230
rect 276 224 282 226
rect 349 226 351 228
rect 353 226 355 228
rect 389 228 395 230
rect 349 224 355 226
rect 389 226 391 228
rect 393 226 395 228
rect 434 228 440 230
rect 389 224 395 226
rect 434 226 436 228
rect 438 226 440 228
rect 434 224 440 226
rect 8 216 14 218
rect 8 214 10 216
rect 12 214 14 216
rect 48 216 54 218
rect 8 212 14 214
rect 48 214 50 216
rect 52 214 54 216
rect 121 216 127 218
rect 48 212 54 214
rect 121 214 123 216
rect 125 214 127 216
rect 152 216 158 218
rect 121 212 127 214
rect 152 214 154 216
rect 156 214 158 216
rect 225 216 231 218
rect 152 212 158 214
rect 225 214 227 216
rect 229 214 231 216
rect 276 216 282 218
rect 225 212 231 214
rect 276 214 278 216
rect 280 214 282 216
rect 349 216 355 218
rect 276 212 282 214
rect 349 214 351 216
rect 353 214 355 216
rect 389 216 395 218
rect 349 212 355 214
rect 389 214 391 216
rect 393 214 395 216
rect 434 216 440 218
rect 389 212 395 214
rect 434 214 436 216
rect 438 214 440 216
rect 434 212 440 214
rect 27 84 33 86
rect 27 82 29 84
rect 31 82 33 84
rect 100 84 106 86
rect 27 80 33 82
rect 100 82 102 84
rect 104 82 106 84
rect 131 84 137 86
rect 100 80 106 82
rect 131 82 133 84
rect 135 82 137 84
rect 204 84 210 86
rect 131 80 137 82
rect 204 82 206 84
rect 208 82 210 84
rect 244 84 250 86
rect 204 80 210 82
rect 244 82 246 84
rect 248 82 250 84
rect 276 84 282 86
rect 244 80 250 82
rect 276 82 278 84
rect 280 82 282 84
rect 349 84 355 86
rect 276 80 282 82
rect 349 82 351 84
rect 353 82 355 84
rect 389 84 395 86
rect 349 80 355 82
rect 389 82 391 84
rect 393 82 395 84
rect 434 84 440 86
rect 389 80 395 82
rect 434 82 436 84
rect 438 82 440 84
rect 434 80 440 82
rect 8 72 14 74
rect 8 70 10 72
rect 12 70 14 72
rect 48 72 54 74
rect 8 68 14 70
rect 48 70 50 72
rect 52 70 54 72
rect 121 72 127 74
rect 48 68 54 70
rect 121 70 123 72
rect 125 70 127 72
rect 152 72 158 74
rect 121 68 127 70
rect 152 70 154 72
rect 156 70 158 72
rect 225 72 231 74
rect 152 68 158 70
rect 225 70 227 72
rect 229 70 231 72
rect 276 72 282 74
rect 225 68 231 70
rect 276 70 278 72
rect 280 70 282 72
rect 349 72 355 74
rect 276 68 282 70
rect 349 70 351 72
rect 353 70 355 72
rect 389 72 395 74
rect 349 68 355 70
rect 389 70 391 72
rect 393 70 395 72
rect 434 72 440 74
rect 389 68 395 70
rect 434 70 436 72
rect 438 70 440 72
rect 434 68 440 70
<< nmos >>
rect 15 560 17 572
rect 22 560 24 572
rect 32 560 34 569
rect 42 560 44 569
rect 58 555 60 564
rect 78 557 80 568
rect 85 557 87 568
rect 98 557 100 566
rect 119 560 121 572
rect 126 560 128 572
rect 136 560 138 569
rect 146 560 148 569
rect 162 555 164 564
rect 182 557 184 568
rect 189 557 191 568
rect 202 557 204 566
rect 222 555 224 561
rect 232 555 234 561
rect 242 555 244 564
rect 264 560 266 572
rect 271 560 273 572
rect 281 560 283 569
rect 291 560 293 569
rect 307 555 309 564
rect 327 557 329 568
rect 334 557 336 568
rect 347 557 349 566
rect 367 555 369 561
rect 377 555 379 561
rect 387 555 389 564
rect 407 555 409 564
rect 423 560 425 569
rect 433 560 435 569
rect 443 560 445 572
rect 450 560 452 572
rect 471 561 473 567
rect 481 561 483 569
rect 488 561 490 569
rect 498 561 500 569
rect 505 561 507 569
rect 515 560 517 569
rect 535 561 537 567
rect 545 561 547 569
rect 552 561 554 569
rect 562 561 564 569
rect 569 561 571 569
rect 579 560 581 569
rect 599 561 601 567
rect 609 561 611 569
rect 616 561 618 569
rect 626 561 628 569
rect 633 561 635 569
rect 643 560 645 569
rect 14 454 16 463
rect 24 457 26 463
rect 34 457 36 463
rect 54 452 56 461
rect 67 450 69 461
rect 74 450 76 461
rect 94 454 96 463
rect 110 449 112 458
rect 120 449 122 458
rect 130 446 132 458
rect 137 446 139 458
rect 158 452 160 461
rect 171 450 173 461
rect 178 450 180 461
rect 198 454 200 463
rect 214 449 216 458
rect 224 449 226 458
rect 234 446 236 458
rect 241 446 243 458
rect 264 446 266 458
rect 271 446 273 458
rect 281 449 283 458
rect 291 449 293 458
rect 307 454 309 463
rect 327 450 329 461
rect 334 450 336 461
rect 347 452 349 461
rect 367 457 369 463
rect 377 457 379 463
rect 387 454 389 463
rect 407 454 409 463
rect 423 449 425 458
rect 433 449 435 458
rect 443 446 445 458
rect 450 446 452 458
rect 471 451 473 457
rect 481 449 483 457
rect 488 449 490 457
rect 498 449 500 457
rect 505 449 507 457
rect 515 449 517 458
rect 535 451 537 457
rect 545 449 547 457
rect 552 449 554 457
rect 562 449 564 457
rect 569 449 571 457
rect 579 449 581 458
rect 599 451 601 457
rect 609 449 611 457
rect 616 449 618 457
rect 626 449 628 457
rect 633 449 635 457
rect 643 449 645 458
rect 15 416 17 428
rect 22 416 24 428
rect 32 416 34 425
rect 42 416 44 425
rect 58 411 60 420
rect 78 413 80 424
rect 85 413 87 424
rect 98 413 100 422
rect 119 416 121 428
rect 126 416 128 428
rect 136 416 138 425
rect 146 416 148 425
rect 162 411 164 420
rect 182 413 184 424
rect 189 413 191 424
rect 202 413 204 422
rect 222 411 224 417
rect 232 411 234 417
rect 242 411 244 420
rect 264 416 266 428
rect 271 416 273 428
rect 281 416 283 425
rect 291 416 293 425
rect 307 411 309 420
rect 327 413 329 424
rect 334 413 336 424
rect 347 413 349 422
rect 367 411 369 417
rect 377 411 379 417
rect 387 411 389 420
rect 407 411 409 420
rect 423 416 425 425
rect 433 416 435 425
rect 443 416 445 428
rect 450 416 452 428
rect 471 417 473 423
rect 481 417 483 425
rect 488 417 490 425
rect 498 417 500 425
rect 505 417 507 425
rect 515 416 517 425
rect 535 417 537 423
rect 545 417 547 425
rect 552 417 554 425
rect 562 417 564 425
rect 569 417 571 425
rect 579 416 581 425
rect 599 417 601 423
rect 609 417 611 425
rect 616 417 618 425
rect 626 417 628 425
rect 633 417 635 425
rect 643 416 645 425
rect 14 310 16 319
rect 24 313 26 319
rect 34 313 36 319
rect 54 308 56 317
rect 67 306 69 317
rect 74 306 76 317
rect 94 310 96 319
rect 110 305 112 314
rect 120 305 122 314
rect 130 302 132 314
rect 137 302 139 314
rect 158 308 160 317
rect 171 306 173 317
rect 178 306 180 317
rect 198 310 200 319
rect 214 305 216 314
rect 224 305 226 314
rect 234 302 236 314
rect 241 302 243 314
rect 264 302 266 314
rect 271 302 273 314
rect 281 305 283 314
rect 291 305 293 314
rect 307 310 309 319
rect 327 306 329 317
rect 334 306 336 317
rect 347 308 349 317
rect 367 313 369 319
rect 377 313 379 319
rect 387 310 389 319
rect 407 310 409 319
rect 423 305 425 314
rect 433 305 435 314
rect 443 302 445 314
rect 450 302 452 314
rect 471 307 473 313
rect 481 305 483 313
rect 488 305 490 313
rect 498 305 500 313
rect 505 305 507 313
rect 515 305 517 314
rect 535 307 537 313
rect 545 305 547 313
rect 552 305 554 313
rect 562 305 564 313
rect 569 305 571 313
rect 579 305 581 314
rect 599 307 601 313
rect 609 305 611 313
rect 616 305 618 313
rect 626 305 628 313
rect 633 305 635 313
rect 643 305 645 314
rect 15 272 17 284
rect 22 272 24 284
rect 32 272 34 281
rect 42 272 44 281
rect 58 267 60 276
rect 78 269 80 280
rect 85 269 87 280
rect 98 269 100 278
rect 119 272 121 284
rect 126 272 128 284
rect 136 272 138 281
rect 146 272 148 281
rect 162 267 164 276
rect 182 269 184 280
rect 189 269 191 280
rect 202 269 204 278
rect 222 267 224 273
rect 232 267 234 273
rect 242 267 244 276
rect 264 272 266 284
rect 271 272 273 284
rect 281 272 283 281
rect 291 272 293 281
rect 307 267 309 276
rect 327 269 329 280
rect 334 269 336 280
rect 347 269 349 278
rect 367 267 369 273
rect 377 267 379 273
rect 387 267 389 276
rect 407 267 409 276
rect 423 272 425 281
rect 433 272 435 281
rect 443 272 445 284
rect 450 272 452 284
rect 471 273 473 279
rect 481 273 483 281
rect 488 273 490 281
rect 498 273 500 281
rect 505 273 507 281
rect 515 272 517 281
rect 535 273 537 279
rect 545 273 547 281
rect 552 273 554 281
rect 562 273 564 281
rect 569 273 571 281
rect 579 272 581 281
rect 599 273 601 279
rect 609 273 611 281
rect 616 273 618 281
rect 626 273 628 281
rect 633 273 635 281
rect 643 272 645 281
rect 14 166 16 175
rect 24 169 26 175
rect 34 169 36 175
rect 54 164 56 173
rect 67 162 69 173
rect 74 162 76 173
rect 94 166 96 175
rect 110 161 112 170
rect 120 161 122 170
rect 130 158 132 170
rect 137 158 139 170
rect 158 164 160 173
rect 171 162 173 173
rect 178 162 180 173
rect 198 166 200 175
rect 214 161 216 170
rect 224 161 226 170
rect 234 158 236 170
rect 241 158 243 170
rect 264 158 266 170
rect 271 158 273 170
rect 281 161 283 170
rect 291 161 293 170
rect 307 166 309 175
rect 327 162 329 173
rect 334 162 336 173
rect 347 164 349 173
rect 367 169 369 175
rect 377 169 379 175
rect 387 166 389 175
rect 407 166 409 175
rect 423 161 425 170
rect 433 161 435 170
rect 443 158 445 170
rect 450 158 452 170
rect 471 163 473 169
rect 481 161 483 169
rect 488 161 490 169
rect 498 161 500 169
rect 505 161 507 169
rect 515 161 517 170
rect 535 163 537 169
rect 545 161 547 169
rect 552 161 554 169
rect 562 161 564 169
rect 569 161 571 169
rect 579 161 581 170
rect 599 163 601 169
rect 609 161 611 169
rect 616 161 618 169
rect 626 161 628 169
rect 633 161 635 169
rect 643 161 645 170
rect 15 128 17 140
rect 22 128 24 140
rect 32 128 34 137
rect 42 128 44 137
rect 58 123 60 132
rect 78 125 80 136
rect 85 125 87 136
rect 98 125 100 134
rect 119 128 121 140
rect 126 128 128 140
rect 136 128 138 137
rect 146 128 148 137
rect 162 123 164 132
rect 182 125 184 136
rect 189 125 191 136
rect 202 125 204 134
rect 222 123 224 129
rect 232 123 234 129
rect 242 123 244 132
rect 264 128 266 140
rect 271 128 273 140
rect 281 128 283 137
rect 291 128 293 137
rect 307 123 309 132
rect 327 125 329 136
rect 334 125 336 136
rect 347 125 349 134
rect 367 123 369 129
rect 377 123 379 129
rect 387 123 389 132
rect 407 123 409 132
rect 423 128 425 137
rect 433 128 435 137
rect 443 128 445 140
rect 450 128 452 140
rect 471 129 473 135
rect 481 129 483 137
rect 488 129 490 137
rect 498 129 500 137
rect 505 129 507 137
rect 515 128 517 137
rect 535 129 537 135
rect 545 129 547 137
rect 552 129 554 137
rect 562 129 564 137
rect 569 129 571 137
rect 579 128 581 137
rect 599 129 601 135
rect 609 129 611 137
rect 616 129 618 137
rect 626 129 628 137
rect 633 129 635 137
rect 643 128 645 137
rect 14 22 16 31
rect 24 25 26 31
rect 34 25 36 31
rect 54 20 56 29
rect 67 18 69 29
rect 74 18 76 29
rect 94 22 96 31
rect 110 17 112 26
rect 120 17 122 26
rect 130 14 132 26
rect 137 14 139 26
rect 158 20 160 29
rect 171 18 173 29
rect 178 18 180 29
rect 198 22 200 31
rect 214 17 216 26
rect 224 17 226 26
rect 234 14 236 26
rect 241 14 243 26
rect 264 14 266 26
rect 271 14 273 26
rect 281 17 283 26
rect 291 17 293 26
rect 307 22 309 31
rect 327 18 329 29
rect 334 18 336 29
rect 347 20 349 29
rect 367 25 369 31
rect 377 25 379 31
rect 387 22 389 31
rect 407 22 409 31
rect 423 17 425 26
rect 433 17 435 26
rect 443 14 445 26
rect 450 14 452 26
rect 471 19 473 25
rect 481 17 483 25
rect 488 17 490 25
rect 498 17 500 25
rect 505 17 507 25
rect 515 17 517 26
rect 535 19 537 25
rect 545 17 547 25
rect 552 17 554 25
rect 562 17 564 25
rect 569 17 571 25
rect 579 17 581 26
rect 599 19 601 25
rect 609 17 611 25
rect 616 17 618 25
rect 626 17 628 25
rect 633 17 635 25
rect 643 17 645 26
<< pmos >>
rect 14 515 16 542
rect 24 524 26 542
rect 34 524 36 542
rect 50 515 52 542
rect 78 522 80 535
rect 88 522 90 535
rect 98 524 100 542
rect 118 515 120 542
rect 128 524 130 542
rect 138 524 140 542
rect 154 515 156 542
rect 182 522 184 535
rect 192 522 194 535
rect 202 524 204 542
rect 222 515 224 536
rect 229 515 231 536
rect 242 525 244 543
rect 263 515 265 542
rect 273 524 275 542
rect 283 524 285 542
rect 299 515 301 542
rect 327 522 329 535
rect 337 522 339 535
rect 347 524 349 542
rect 367 515 369 536
rect 374 515 376 536
rect 387 525 389 543
rect 415 515 417 542
rect 431 524 433 542
rect 441 524 443 542
rect 451 515 453 542
rect 471 535 473 543
rect 535 535 537 543
rect 481 515 483 531
rect 488 515 490 531
rect 498 515 500 531
rect 505 515 507 531
rect 515 515 517 533
rect 599 535 601 543
rect 545 515 547 531
rect 552 515 554 531
rect 562 515 564 531
rect 569 515 571 531
rect 579 515 581 533
rect 609 515 611 531
rect 616 515 618 531
rect 626 515 628 531
rect 633 515 635 531
rect 643 515 645 533
rect 14 475 16 493
rect 27 482 29 503
rect 34 482 36 503
rect 54 476 56 494
rect 64 483 66 496
rect 74 483 76 496
rect 102 476 104 503
rect 118 476 120 494
rect 128 476 130 494
rect 138 476 140 503
rect 158 476 160 494
rect 168 483 170 496
rect 178 483 180 496
rect 206 476 208 503
rect 222 476 224 494
rect 232 476 234 494
rect 242 476 244 503
rect 263 476 265 503
rect 273 476 275 494
rect 283 476 285 494
rect 299 476 301 503
rect 327 483 329 496
rect 337 483 339 496
rect 347 476 349 494
rect 367 482 369 503
rect 374 482 376 503
rect 387 475 389 493
rect 415 476 417 503
rect 431 476 433 494
rect 441 476 443 494
rect 451 476 453 503
rect 481 487 483 503
rect 488 487 490 503
rect 498 487 500 503
rect 505 487 507 503
rect 471 475 473 483
rect 515 485 517 503
rect 545 487 547 503
rect 552 487 554 503
rect 562 487 564 503
rect 569 487 571 503
rect 535 475 537 483
rect 579 485 581 503
rect 609 487 611 503
rect 616 487 618 503
rect 626 487 628 503
rect 633 487 635 503
rect 599 475 601 483
rect 643 485 645 503
rect 14 371 16 398
rect 24 380 26 398
rect 34 380 36 398
rect 50 371 52 398
rect 78 378 80 391
rect 88 378 90 391
rect 98 380 100 398
rect 118 371 120 398
rect 128 380 130 398
rect 138 380 140 398
rect 154 371 156 398
rect 182 378 184 391
rect 192 378 194 391
rect 202 380 204 398
rect 222 371 224 392
rect 229 371 231 392
rect 242 381 244 399
rect 263 371 265 398
rect 273 380 275 398
rect 283 380 285 398
rect 299 371 301 398
rect 327 378 329 391
rect 337 378 339 391
rect 347 380 349 398
rect 367 371 369 392
rect 374 371 376 392
rect 387 381 389 399
rect 415 371 417 398
rect 431 380 433 398
rect 441 380 443 398
rect 451 371 453 398
rect 471 391 473 399
rect 535 391 537 399
rect 481 371 483 387
rect 488 371 490 387
rect 498 371 500 387
rect 505 371 507 387
rect 515 371 517 389
rect 599 391 601 399
rect 545 371 547 387
rect 552 371 554 387
rect 562 371 564 387
rect 569 371 571 387
rect 579 371 581 389
rect 609 371 611 387
rect 616 371 618 387
rect 626 371 628 387
rect 633 371 635 387
rect 643 371 645 389
rect 14 331 16 349
rect 27 338 29 359
rect 34 338 36 359
rect 54 332 56 350
rect 64 339 66 352
rect 74 339 76 352
rect 102 332 104 359
rect 118 332 120 350
rect 128 332 130 350
rect 138 332 140 359
rect 158 332 160 350
rect 168 339 170 352
rect 178 339 180 352
rect 206 332 208 359
rect 222 332 224 350
rect 232 332 234 350
rect 242 332 244 359
rect 263 332 265 359
rect 273 332 275 350
rect 283 332 285 350
rect 299 332 301 359
rect 327 339 329 352
rect 337 339 339 352
rect 347 332 349 350
rect 367 338 369 359
rect 374 338 376 359
rect 387 331 389 349
rect 415 332 417 359
rect 431 332 433 350
rect 441 332 443 350
rect 451 332 453 359
rect 481 343 483 359
rect 488 343 490 359
rect 498 343 500 359
rect 505 343 507 359
rect 471 331 473 339
rect 515 341 517 359
rect 545 343 547 359
rect 552 343 554 359
rect 562 343 564 359
rect 569 343 571 359
rect 535 331 537 339
rect 579 341 581 359
rect 609 343 611 359
rect 616 343 618 359
rect 626 343 628 359
rect 633 343 635 359
rect 599 331 601 339
rect 643 341 645 359
rect 14 227 16 254
rect 24 236 26 254
rect 34 236 36 254
rect 50 227 52 254
rect 78 234 80 247
rect 88 234 90 247
rect 98 236 100 254
rect 118 227 120 254
rect 128 236 130 254
rect 138 236 140 254
rect 154 227 156 254
rect 182 234 184 247
rect 192 234 194 247
rect 202 236 204 254
rect 222 227 224 248
rect 229 227 231 248
rect 242 237 244 255
rect 263 227 265 254
rect 273 236 275 254
rect 283 236 285 254
rect 299 227 301 254
rect 327 234 329 247
rect 337 234 339 247
rect 347 236 349 254
rect 367 227 369 248
rect 374 227 376 248
rect 387 237 389 255
rect 415 227 417 254
rect 431 236 433 254
rect 441 236 443 254
rect 451 227 453 254
rect 471 247 473 255
rect 535 247 537 255
rect 481 227 483 243
rect 488 227 490 243
rect 498 227 500 243
rect 505 227 507 243
rect 515 227 517 245
rect 599 247 601 255
rect 545 227 547 243
rect 552 227 554 243
rect 562 227 564 243
rect 569 227 571 243
rect 579 227 581 245
rect 609 227 611 243
rect 616 227 618 243
rect 626 227 628 243
rect 633 227 635 243
rect 643 227 645 245
rect 14 187 16 205
rect 27 194 29 215
rect 34 194 36 215
rect 54 188 56 206
rect 64 195 66 208
rect 74 195 76 208
rect 102 188 104 215
rect 118 188 120 206
rect 128 188 130 206
rect 138 188 140 215
rect 158 188 160 206
rect 168 195 170 208
rect 178 195 180 208
rect 206 188 208 215
rect 222 188 224 206
rect 232 188 234 206
rect 242 188 244 215
rect 263 188 265 215
rect 273 188 275 206
rect 283 188 285 206
rect 299 188 301 215
rect 327 195 329 208
rect 337 195 339 208
rect 347 188 349 206
rect 367 194 369 215
rect 374 194 376 215
rect 387 187 389 205
rect 415 188 417 215
rect 431 188 433 206
rect 441 188 443 206
rect 451 188 453 215
rect 481 199 483 215
rect 488 199 490 215
rect 498 199 500 215
rect 505 199 507 215
rect 471 187 473 195
rect 515 197 517 215
rect 545 199 547 215
rect 552 199 554 215
rect 562 199 564 215
rect 569 199 571 215
rect 535 187 537 195
rect 579 197 581 215
rect 609 199 611 215
rect 616 199 618 215
rect 626 199 628 215
rect 633 199 635 215
rect 599 187 601 195
rect 643 197 645 215
rect 14 83 16 110
rect 24 92 26 110
rect 34 92 36 110
rect 50 83 52 110
rect 78 90 80 103
rect 88 90 90 103
rect 98 92 100 110
rect 118 83 120 110
rect 128 92 130 110
rect 138 92 140 110
rect 154 83 156 110
rect 182 90 184 103
rect 192 90 194 103
rect 202 92 204 110
rect 222 83 224 104
rect 229 83 231 104
rect 242 93 244 111
rect 263 83 265 110
rect 273 92 275 110
rect 283 92 285 110
rect 299 83 301 110
rect 327 90 329 103
rect 337 90 339 103
rect 347 92 349 110
rect 367 83 369 104
rect 374 83 376 104
rect 387 93 389 111
rect 415 83 417 110
rect 431 92 433 110
rect 441 92 443 110
rect 451 83 453 110
rect 471 103 473 111
rect 535 103 537 111
rect 481 83 483 99
rect 488 83 490 99
rect 498 83 500 99
rect 505 83 507 99
rect 515 83 517 101
rect 599 103 601 111
rect 545 83 547 99
rect 552 83 554 99
rect 562 83 564 99
rect 569 83 571 99
rect 579 83 581 101
rect 609 83 611 99
rect 616 83 618 99
rect 626 83 628 99
rect 633 83 635 99
rect 643 83 645 101
rect 14 43 16 61
rect 27 50 29 71
rect 34 50 36 71
rect 54 44 56 62
rect 64 51 66 64
rect 74 51 76 64
rect 102 44 104 71
rect 118 44 120 62
rect 128 44 130 62
rect 138 44 140 71
rect 158 44 160 62
rect 168 51 170 64
rect 178 51 180 64
rect 206 44 208 71
rect 222 44 224 62
rect 232 44 234 62
rect 242 44 244 71
rect 263 44 265 71
rect 273 44 275 62
rect 283 44 285 62
rect 299 44 301 71
rect 327 51 329 64
rect 337 51 339 64
rect 347 44 349 62
rect 367 50 369 71
rect 374 50 376 71
rect 387 43 389 61
rect 415 44 417 71
rect 431 44 433 62
rect 441 44 443 62
rect 451 44 453 71
rect 481 55 483 71
rect 488 55 490 71
rect 498 55 500 71
rect 505 55 507 71
rect 471 43 473 51
rect 515 53 517 71
rect 545 55 547 71
rect 552 55 554 71
rect 562 55 564 71
rect 569 55 571 71
rect 535 43 537 51
rect 579 53 581 71
rect 609 55 611 71
rect 616 55 618 71
rect 626 55 628 71
rect 633 55 635 71
rect 599 43 601 51
rect 643 53 645 71
<< polyct0 >>
rect 16 547 18 549
rect 26 548 28 550
rect 96 548 98 550
rect 120 547 122 549
rect 130 548 132 550
rect 200 548 202 550
rect 240 548 242 550
rect 265 547 267 549
rect 275 548 277 550
rect 345 548 347 550
rect 385 548 387 550
rect 439 548 441 550
rect 449 547 451 549
rect 496 554 498 556
rect 514 553 516 555
rect 489 538 491 540
rect 560 554 562 556
rect 578 553 580 555
rect 553 538 555 540
rect 624 554 626 556
rect 642 553 644 555
rect 617 538 619 540
rect 16 468 18 470
rect 56 468 58 470
rect 126 468 128 470
rect 136 469 138 471
rect 160 468 162 470
rect 230 468 232 470
rect 240 469 242 471
rect 265 469 267 471
rect 275 468 277 470
rect 345 468 347 470
rect 385 468 387 470
rect 439 468 441 470
rect 449 469 451 471
rect 489 478 491 480
rect 496 462 498 464
rect 514 463 516 465
rect 553 478 555 480
rect 560 462 562 464
rect 578 463 580 465
rect 617 478 619 480
rect 624 462 626 464
rect 642 463 644 465
rect 16 403 18 405
rect 26 404 28 406
rect 96 404 98 406
rect 120 403 122 405
rect 130 404 132 406
rect 200 404 202 406
rect 240 404 242 406
rect 265 403 267 405
rect 275 404 277 406
rect 345 404 347 406
rect 385 404 387 406
rect 439 404 441 406
rect 449 403 451 405
rect 496 410 498 412
rect 514 409 516 411
rect 489 394 491 396
rect 560 410 562 412
rect 578 409 580 411
rect 553 394 555 396
rect 624 410 626 412
rect 642 409 644 411
rect 617 394 619 396
rect 16 324 18 326
rect 56 324 58 326
rect 126 324 128 326
rect 136 325 138 327
rect 160 324 162 326
rect 230 324 232 326
rect 240 325 242 327
rect 265 325 267 327
rect 275 324 277 326
rect 345 324 347 326
rect 385 324 387 326
rect 439 324 441 326
rect 449 325 451 327
rect 489 334 491 336
rect 496 318 498 320
rect 514 319 516 321
rect 553 334 555 336
rect 560 318 562 320
rect 578 319 580 321
rect 617 334 619 336
rect 624 318 626 320
rect 642 319 644 321
rect 16 259 18 261
rect 26 260 28 262
rect 96 260 98 262
rect 120 259 122 261
rect 130 260 132 262
rect 200 260 202 262
rect 240 260 242 262
rect 265 259 267 261
rect 275 260 277 262
rect 345 260 347 262
rect 385 260 387 262
rect 439 260 441 262
rect 449 259 451 261
rect 496 266 498 268
rect 514 265 516 267
rect 489 250 491 252
rect 560 266 562 268
rect 578 265 580 267
rect 553 250 555 252
rect 624 266 626 268
rect 642 265 644 267
rect 617 250 619 252
rect 16 180 18 182
rect 56 180 58 182
rect 126 180 128 182
rect 136 181 138 183
rect 160 180 162 182
rect 230 180 232 182
rect 240 181 242 183
rect 265 181 267 183
rect 275 180 277 182
rect 345 180 347 182
rect 385 180 387 182
rect 439 180 441 182
rect 449 181 451 183
rect 489 190 491 192
rect 496 174 498 176
rect 514 175 516 177
rect 553 190 555 192
rect 560 174 562 176
rect 578 175 580 177
rect 617 190 619 192
rect 624 174 626 176
rect 642 175 644 177
rect 16 115 18 117
rect 26 116 28 118
rect 96 116 98 118
rect 120 115 122 117
rect 130 116 132 118
rect 200 116 202 118
rect 240 116 242 118
rect 265 115 267 117
rect 275 116 277 118
rect 345 116 347 118
rect 385 116 387 118
rect 439 116 441 118
rect 449 115 451 117
rect 496 122 498 124
rect 514 121 516 123
rect 489 106 491 108
rect 560 122 562 124
rect 578 121 580 123
rect 553 106 555 108
rect 624 122 626 124
rect 642 121 644 123
rect 617 106 619 108
rect 16 36 18 38
rect 56 36 58 38
rect 126 36 128 38
rect 136 37 138 39
rect 160 36 162 38
rect 230 36 232 38
rect 240 37 242 39
rect 265 37 267 39
rect 275 36 277 38
rect 345 36 347 38
rect 385 36 387 38
rect 439 36 441 38
rect 449 37 451 39
rect 489 46 491 48
rect 496 30 498 32
rect 514 31 516 33
rect 553 46 555 48
rect 560 30 562 32
rect 578 31 580 33
rect 617 46 619 48
rect 624 30 626 32
rect 642 31 644 33
<< polyct1 >>
rect 47 553 49 555
rect 86 548 88 550
rect 151 553 153 555
rect 63 540 65 542
rect 76 540 78 542
rect 190 548 192 550
rect 167 540 169 542
rect 180 540 182 542
rect 230 548 232 550
rect 296 553 298 555
rect 220 541 222 543
rect 335 548 337 550
rect 312 540 314 542
rect 325 540 327 542
rect 375 548 377 550
rect 418 553 420 555
rect 365 541 367 543
rect 479 548 481 550
rect 402 540 404 542
rect 506 543 508 545
rect 543 548 545 550
rect 466 528 468 530
rect 570 543 572 545
rect 607 548 609 550
rect 530 528 532 530
rect 634 543 636 545
rect 594 528 596 530
rect 36 475 38 477
rect 26 468 28 470
rect 76 476 78 478
rect 89 476 91 478
rect 66 468 68 470
rect 180 476 182 478
rect 193 476 195 478
rect 312 476 314 478
rect 105 463 107 465
rect 170 468 172 470
rect 325 476 327 478
rect 209 463 211 465
rect 296 463 298 465
rect 365 475 367 477
rect 335 468 337 470
rect 402 476 404 478
rect 466 488 468 490
rect 375 468 377 470
rect 418 463 420 465
rect 530 488 532 490
rect 479 468 481 470
rect 506 473 508 475
rect 594 488 596 490
rect 543 468 545 470
rect 570 473 572 475
rect 607 468 609 470
rect 634 473 636 475
rect 47 409 49 411
rect 86 404 88 406
rect 151 409 153 411
rect 63 396 65 398
rect 76 396 78 398
rect 190 404 192 406
rect 167 396 169 398
rect 180 396 182 398
rect 230 404 232 406
rect 296 409 298 411
rect 220 397 222 399
rect 335 404 337 406
rect 312 396 314 398
rect 325 396 327 398
rect 375 404 377 406
rect 418 409 420 411
rect 365 397 367 399
rect 479 404 481 406
rect 402 396 404 398
rect 506 399 508 401
rect 543 404 545 406
rect 466 384 468 386
rect 570 399 572 401
rect 607 404 609 406
rect 530 384 532 386
rect 634 399 636 401
rect 594 384 596 386
rect 36 331 38 333
rect 26 324 28 326
rect 76 332 78 334
rect 89 332 91 334
rect 66 324 68 326
rect 180 332 182 334
rect 193 332 195 334
rect 312 332 314 334
rect 105 319 107 321
rect 170 324 172 326
rect 325 332 327 334
rect 209 319 211 321
rect 296 319 298 321
rect 365 331 367 333
rect 335 324 337 326
rect 402 332 404 334
rect 466 344 468 346
rect 375 324 377 326
rect 418 319 420 321
rect 530 344 532 346
rect 479 324 481 326
rect 506 329 508 331
rect 594 344 596 346
rect 543 324 545 326
rect 570 329 572 331
rect 607 324 609 326
rect 634 329 636 331
rect 47 265 49 267
rect 86 260 88 262
rect 151 265 153 267
rect 63 252 65 254
rect 76 252 78 254
rect 190 260 192 262
rect 167 252 169 254
rect 180 252 182 254
rect 230 260 232 262
rect 296 265 298 267
rect 220 253 222 255
rect 335 260 337 262
rect 312 252 314 254
rect 325 252 327 254
rect 375 260 377 262
rect 418 265 420 267
rect 365 253 367 255
rect 479 260 481 262
rect 402 252 404 254
rect 506 255 508 257
rect 543 260 545 262
rect 466 240 468 242
rect 570 255 572 257
rect 607 260 609 262
rect 530 240 532 242
rect 634 255 636 257
rect 594 240 596 242
rect 36 187 38 189
rect 26 180 28 182
rect 76 188 78 190
rect 89 188 91 190
rect 66 180 68 182
rect 180 188 182 190
rect 193 188 195 190
rect 312 188 314 190
rect 105 175 107 177
rect 170 180 172 182
rect 325 188 327 190
rect 209 175 211 177
rect 296 175 298 177
rect 365 187 367 189
rect 335 180 337 182
rect 402 188 404 190
rect 466 200 468 202
rect 375 180 377 182
rect 418 175 420 177
rect 530 200 532 202
rect 479 180 481 182
rect 506 185 508 187
rect 594 200 596 202
rect 543 180 545 182
rect 570 185 572 187
rect 607 180 609 182
rect 634 185 636 187
rect 47 121 49 123
rect 86 116 88 118
rect 151 121 153 123
rect 63 108 65 110
rect 76 108 78 110
rect 190 116 192 118
rect 167 108 169 110
rect 180 108 182 110
rect 230 116 232 118
rect 296 121 298 123
rect 220 109 222 111
rect 335 116 337 118
rect 312 108 314 110
rect 325 108 327 110
rect 375 116 377 118
rect 418 121 420 123
rect 365 109 367 111
rect 479 116 481 118
rect 402 108 404 110
rect 506 111 508 113
rect 543 116 545 118
rect 466 96 468 98
rect 570 111 572 113
rect 607 116 609 118
rect 530 96 532 98
rect 634 111 636 113
rect 594 96 596 98
rect 36 43 38 45
rect 26 36 28 38
rect 76 44 78 46
rect 89 44 91 46
rect 66 36 68 38
rect 180 44 182 46
rect 193 44 195 46
rect 312 44 314 46
rect 105 31 107 33
rect 170 36 172 38
rect 325 44 327 46
rect 209 31 211 33
rect 296 31 298 33
rect 365 43 367 45
rect 335 36 337 38
rect 402 44 404 46
rect 466 56 468 58
rect 375 36 377 38
rect 418 31 420 33
rect 530 56 532 58
rect 479 36 481 38
rect 506 41 508 43
rect 594 56 596 58
rect 543 36 545 38
rect 570 41 572 43
rect 607 36 609 38
rect 634 41 636 43
<< ndifct0 >>
rect 37 562 39 564
rect 49 565 51 567
rect 73 564 75 566
rect 63 557 65 559
rect 141 562 143 564
rect 217 570 219 572
rect 153 565 155 567
rect 177 564 179 566
rect 167 557 169 559
rect 236 570 238 572
rect 227 557 229 559
rect 286 562 288 564
rect 362 570 364 572
rect 298 565 300 567
rect 322 564 324 566
rect 312 557 314 559
rect 381 570 383 572
rect 416 565 418 567
rect 372 557 374 559
rect 402 557 404 559
rect 428 562 430 564
rect 466 563 468 565
rect 476 563 478 565
rect 493 565 495 567
rect 510 565 512 567
rect 530 563 532 565
rect 540 563 542 565
rect 557 565 559 567
rect 574 565 576 567
rect 594 563 596 565
rect 604 563 606 565
rect 621 565 623 567
rect 638 565 640 567
rect 29 459 31 461
rect 20 446 22 448
rect 89 459 91 461
rect 79 452 81 454
rect 103 451 105 453
rect 39 446 41 448
rect 115 454 117 456
rect 193 459 195 461
rect 183 452 185 454
rect 207 451 209 453
rect 219 454 221 456
rect 286 454 288 456
rect 312 459 314 461
rect 298 451 300 453
rect 322 452 324 454
rect 372 459 374 461
rect 402 459 404 461
rect 362 446 364 448
rect 416 451 418 453
rect 428 454 430 456
rect 381 446 383 448
rect 466 453 468 455
rect 476 453 478 455
rect 493 451 495 453
rect 510 451 512 453
rect 530 453 532 455
rect 540 453 542 455
rect 557 451 559 453
rect 574 451 576 453
rect 594 453 596 455
rect 604 453 606 455
rect 621 451 623 453
rect 638 451 640 453
rect 37 418 39 420
rect 49 421 51 423
rect 73 420 75 422
rect 63 413 65 415
rect 141 418 143 420
rect 217 426 219 428
rect 153 421 155 423
rect 177 420 179 422
rect 167 413 169 415
rect 236 426 238 428
rect 227 413 229 415
rect 286 418 288 420
rect 362 426 364 428
rect 298 421 300 423
rect 322 420 324 422
rect 312 413 314 415
rect 381 426 383 428
rect 416 421 418 423
rect 372 413 374 415
rect 402 413 404 415
rect 428 418 430 420
rect 466 419 468 421
rect 476 419 478 421
rect 493 421 495 423
rect 510 421 512 423
rect 530 419 532 421
rect 540 419 542 421
rect 557 421 559 423
rect 574 421 576 423
rect 594 419 596 421
rect 604 419 606 421
rect 621 421 623 423
rect 638 421 640 423
rect 29 315 31 317
rect 20 302 22 304
rect 89 315 91 317
rect 79 308 81 310
rect 103 307 105 309
rect 39 302 41 304
rect 115 310 117 312
rect 193 315 195 317
rect 183 308 185 310
rect 207 307 209 309
rect 219 310 221 312
rect 286 310 288 312
rect 312 315 314 317
rect 298 307 300 309
rect 322 308 324 310
rect 372 315 374 317
rect 402 315 404 317
rect 362 302 364 304
rect 416 307 418 309
rect 428 310 430 312
rect 381 302 383 304
rect 466 309 468 311
rect 476 309 478 311
rect 493 307 495 309
rect 510 307 512 309
rect 530 309 532 311
rect 540 309 542 311
rect 557 307 559 309
rect 574 307 576 309
rect 594 309 596 311
rect 604 309 606 311
rect 621 307 623 309
rect 638 307 640 309
rect 37 274 39 276
rect 49 277 51 279
rect 73 276 75 278
rect 63 269 65 271
rect 141 274 143 276
rect 217 282 219 284
rect 153 277 155 279
rect 177 276 179 278
rect 167 269 169 271
rect 236 282 238 284
rect 227 269 229 271
rect 286 274 288 276
rect 362 282 364 284
rect 298 277 300 279
rect 322 276 324 278
rect 312 269 314 271
rect 381 282 383 284
rect 416 277 418 279
rect 372 269 374 271
rect 402 269 404 271
rect 428 274 430 276
rect 466 275 468 277
rect 476 275 478 277
rect 493 277 495 279
rect 510 277 512 279
rect 530 275 532 277
rect 540 275 542 277
rect 557 277 559 279
rect 574 277 576 279
rect 594 275 596 277
rect 604 275 606 277
rect 621 277 623 279
rect 638 277 640 279
rect 29 171 31 173
rect 20 158 22 160
rect 89 171 91 173
rect 79 164 81 166
rect 103 163 105 165
rect 39 158 41 160
rect 115 166 117 168
rect 193 171 195 173
rect 183 164 185 166
rect 207 163 209 165
rect 219 166 221 168
rect 286 166 288 168
rect 312 171 314 173
rect 298 163 300 165
rect 322 164 324 166
rect 372 171 374 173
rect 402 171 404 173
rect 362 158 364 160
rect 416 163 418 165
rect 428 166 430 168
rect 381 158 383 160
rect 466 165 468 167
rect 476 165 478 167
rect 493 163 495 165
rect 510 163 512 165
rect 530 165 532 167
rect 540 165 542 167
rect 557 163 559 165
rect 574 163 576 165
rect 594 165 596 167
rect 604 165 606 167
rect 621 163 623 165
rect 638 163 640 165
rect 37 130 39 132
rect 49 133 51 135
rect 73 132 75 134
rect 63 125 65 127
rect 141 130 143 132
rect 217 138 219 140
rect 153 133 155 135
rect 177 132 179 134
rect 167 125 169 127
rect 236 138 238 140
rect 227 125 229 127
rect 286 130 288 132
rect 362 138 364 140
rect 298 133 300 135
rect 322 132 324 134
rect 312 125 314 127
rect 381 138 383 140
rect 416 133 418 135
rect 372 125 374 127
rect 402 125 404 127
rect 428 130 430 132
rect 466 131 468 133
rect 476 131 478 133
rect 493 133 495 135
rect 510 133 512 135
rect 530 131 532 133
rect 540 131 542 133
rect 557 133 559 135
rect 574 133 576 135
rect 594 131 596 133
rect 604 131 606 133
rect 621 133 623 135
rect 638 133 640 135
rect 29 27 31 29
rect 20 14 22 16
rect 89 27 91 29
rect 79 20 81 22
rect 103 19 105 21
rect 39 14 41 16
rect 115 22 117 24
rect 193 27 195 29
rect 183 20 185 22
rect 207 19 209 21
rect 219 22 221 24
rect 286 22 288 24
rect 312 27 314 29
rect 298 19 300 21
rect 322 20 324 22
rect 372 27 374 29
rect 402 27 404 29
rect 362 14 364 16
rect 416 19 418 21
rect 428 22 430 24
rect 381 14 383 16
rect 466 21 468 23
rect 476 21 478 23
rect 493 19 495 21
rect 510 19 512 21
rect 530 21 532 23
rect 540 21 542 23
rect 557 19 559 21
rect 574 19 576 21
rect 594 21 596 23
rect 604 21 606 23
rect 621 19 623 21
rect 638 19 640 21
<< ndifct1 >>
rect 9 574 11 576
rect 92 574 94 576
rect 27 564 29 566
rect 113 574 115 576
rect 103 562 105 564
rect 196 574 198 576
rect 131 564 133 566
rect 258 574 260 576
rect 207 562 209 564
rect 341 574 343 576
rect 276 564 278 566
rect 247 557 249 559
rect 456 574 458 576
rect 352 562 354 564
rect 392 557 394 559
rect 438 564 440 566
rect 520 562 522 564
rect 584 562 586 564
rect 648 562 650 564
rect 9 459 11 461
rect 49 454 51 456
rect 125 452 127 454
rect 60 442 62 444
rect 153 454 155 456
rect 143 442 145 444
rect 229 452 231 454
rect 164 442 166 444
rect 247 442 249 444
rect 276 452 278 454
rect 352 454 354 456
rect 258 442 260 444
rect 392 459 394 461
rect 341 442 343 444
rect 438 452 440 454
rect 456 442 458 444
rect 520 454 522 456
rect 584 454 586 456
rect 648 454 650 456
rect 9 430 11 432
rect 92 430 94 432
rect 27 420 29 422
rect 113 430 115 432
rect 103 418 105 420
rect 196 430 198 432
rect 131 420 133 422
rect 258 430 260 432
rect 207 418 209 420
rect 341 430 343 432
rect 276 420 278 422
rect 247 413 249 415
rect 456 430 458 432
rect 352 418 354 420
rect 392 413 394 415
rect 438 420 440 422
rect 520 418 522 420
rect 584 418 586 420
rect 648 418 650 420
rect 9 315 11 317
rect 49 310 51 312
rect 125 308 127 310
rect 60 298 62 300
rect 153 310 155 312
rect 143 298 145 300
rect 229 308 231 310
rect 164 298 166 300
rect 247 298 249 300
rect 276 308 278 310
rect 352 310 354 312
rect 258 298 260 300
rect 392 315 394 317
rect 341 298 343 300
rect 438 308 440 310
rect 456 298 458 300
rect 520 310 522 312
rect 584 310 586 312
rect 648 310 650 312
rect 9 286 11 288
rect 92 286 94 288
rect 27 276 29 278
rect 113 286 115 288
rect 103 274 105 276
rect 196 286 198 288
rect 131 276 133 278
rect 258 286 260 288
rect 207 274 209 276
rect 341 286 343 288
rect 276 276 278 278
rect 247 269 249 271
rect 456 286 458 288
rect 352 274 354 276
rect 392 269 394 271
rect 438 276 440 278
rect 520 274 522 276
rect 584 274 586 276
rect 648 274 650 276
rect 9 171 11 173
rect 49 166 51 168
rect 125 164 127 166
rect 60 154 62 156
rect 153 166 155 168
rect 143 154 145 156
rect 229 164 231 166
rect 164 154 166 156
rect 247 154 249 156
rect 276 164 278 166
rect 352 166 354 168
rect 258 154 260 156
rect 392 171 394 173
rect 341 154 343 156
rect 438 164 440 166
rect 456 154 458 156
rect 520 166 522 168
rect 584 166 586 168
rect 648 166 650 168
rect 9 142 11 144
rect 92 142 94 144
rect 27 132 29 134
rect 113 142 115 144
rect 103 130 105 132
rect 196 142 198 144
rect 131 132 133 134
rect 258 142 260 144
rect 207 130 209 132
rect 341 142 343 144
rect 276 132 278 134
rect 247 125 249 127
rect 456 142 458 144
rect 352 130 354 132
rect 392 125 394 127
rect 438 132 440 134
rect 520 130 522 132
rect 584 130 586 132
rect 648 130 650 132
rect 9 27 11 29
rect 49 22 51 24
rect 125 20 127 22
rect 60 10 62 12
rect 153 22 155 24
rect 143 10 145 12
rect 229 20 231 22
rect 164 10 166 12
rect 247 10 249 12
rect 276 20 278 22
rect 352 22 354 24
rect 258 10 260 12
rect 392 27 394 29
rect 341 10 343 12
rect 438 20 440 22
rect 456 10 458 12
rect 520 22 522 24
rect 584 22 586 24
rect 648 22 650 24
<< ntiect1 >>
rect 29 514 31 516
rect 102 514 104 516
rect 133 514 135 516
rect 206 514 208 516
rect 246 514 248 516
rect 278 514 280 516
rect 351 514 353 516
rect 391 514 393 516
rect 436 514 438 516
rect 10 502 12 504
rect 50 502 52 504
rect 123 502 125 504
rect 154 502 156 504
rect 227 502 229 504
rect 278 502 280 504
rect 351 502 353 504
rect 391 502 393 504
rect 436 502 438 504
rect 29 370 31 372
rect 102 370 104 372
rect 133 370 135 372
rect 206 370 208 372
rect 246 370 248 372
rect 278 370 280 372
rect 351 370 353 372
rect 391 370 393 372
rect 436 370 438 372
rect 10 358 12 360
rect 50 358 52 360
rect 123 358 125 360
rect 154 358 156 360
rect 227 358 229 360
rect 278 358 280 360
rect 351 358 353 360
rect 391 358 393 360
rect 436 358 438 360
rect 29 226 31 228
rect 102 226 104 228
rect 133 226 135 228
rect 206 226 208 228
rect 246 226 248 228
rect 278 226 280 228
rect 351 226 353 228
rect 391 226 393 228
rect 436 226 438 228
rect 10 214 12 216
rect 50 214 52 216
rect 123 214 125 216
rect 154 214 156 216
rect 227 214 229 216
rect 278 214 280 216
rect 351 214 353 216
rect 391 214 393 216
rect 436 214 438 216
rect 29 82 31 84
rect 102 82 104 84
rect 133 82 135 84
rect 206 82 208 84
rect 246 82 248 84
rect 278 82 280 84
rect 351 82 353 84
rect 391 82 393 84
rect 436 82 438 84
rect 10 70 12 72
rect 50 70 52 72
rect 123 70 125 72
rect 154 70 156 72
rect 227 70 229 72
rect 278 70 280 72
rect 351 70 353 72
rect 391 70 393 72
rect 436 70 438 72
<< ptiect1 >>
rect 62 574 64 576
rect 102 574 104 576
rect 166 574 168 576
rect 206 574 208 576
rect 246 574 248 576
rect 311 574 313 576
rect 351 574 353 576
rect 391 574 393 576
rect 403 574 405 576
rect 10 442 12 444
rect 50 442 52 444
rect 90 442 92 444
rect 154 442 156 444
rect 194 442 196 444
rect 311 442 313 444
rect 351 442 353 444
rect 391 442 393 444
rect 403 442 405 444
rect 62 430 64 432
rect 102 430 104 432
rect 166 430 168 432
rect 206 430 208 432
rect 246 430 248 432
rect 311 430 313 432
rect 351 430 353 432
rect 391 430 393 432
rect 403 430 405 432
rect 10 298 12 300
rect 50 298 52 300
rect 90 298 92 300
rect 154 298 156 300
rect 194 298 196 300
rect 311 298 313 300
rect 351 298 353 300
rect 391 298 393 300
rect 403 298 405 300
rect 62 286 64 288
rect 102 286 104 288
rect 166 286 168 288
rect 206 286 208 288
rect 246 286 248 288
rect 311 286 313 288
rect 351 286 353 288
rect 391 286 393 288
rect 403 286 405 288
rect 10 154 12 156
rect 50 154 52 156
rect 90 154 92 156
rect 154 154 156 156
rect 194 154 196 156
rect 311 154 313 156
rect 351 154 353 156
rect 391 154 393 156
rect 403 154 405 156
rect 62 142 64 144
rect 102 142 104 144
rect 166 142 168 144
rect 206 142 208 144
rect 246 142 248 144
rect 311 142 313 144
rect 351 142 353 144
rect 391 142 393 144
rect 403 142 405 144
rect 10 10 12 12
rect 50 10 52 12
rect 90 10 92 12
rect 154 10 156 12
rect 194 10 196 12
rect 311 10 313 12
rect 351 10 353 12
rect 391 10 393 12
rect 403 10 405 12
<< pdifct0 >>
rect 9 523 11 525
rect 29 538 31 540
rect 29 531 31 533
rect 45 524 47 526
rect 45 517 47 519
rect 55 538 57 540
rect 73 524 75 526
rect 83 531 85 533
rect 83 524 85 526
rect 93 526 95 528
rect 113 523 115 525
rect 133 538 135 540
rect 133 531 135 533
rect 149 524 151 526
rect 149 517 151 519
rect 159 538 161 540
rect 177 524 179 526
rect 187 531 189 533
rect 187 524 189 526
rect 197 526 199 528
rect 217 524 219 526
rect 258 523 260 525
rect 236 517 238 519
rect 278 538 280 540
rect 278 531 280 533
rect 294 524 296 526
rect 294 517 296 519
rect 304 538 306 540
rect 322 524 324 526
rect 332 531 334 533
rect 332 524 334 526
rect 342 526 344 528
rect 362 524 364 526
rect 410 538 412 540
rect 381 517 383 519
rect 420 524 422 526
rect 436 538 438 540
rect 436 531 438 533
rect 420 517 422 519
rect 466 539 468 541
rect 530 539 532 541
rect 456 523 458 525
rect 476 517 478 519
rect 493 527 495 529
rect 510 517 512 519
rect 594 539 596 541
rect 540 517 542 519
rect 557 527 559 529
rect 574 517 576 519
rect 604 517 606 519
rect 621 527 623 529
rect 638 517 640 519
rect 20 499 22 501
rect 39 492 41 494
rect 59 490 61 492
rect 69 492 71 494
rect 69 485 71 487
rect 79 492 81 494
rect 97 478 99 480
rect 107 499 109 501
rect 107 492 109 494
rect 123 485 125 487
rect 123 478 125 480
rect 143 493 145 495
rect 163 490 165 492
rect 173 492 175 494
rect 173 485 175 487
rect 183 492 185 494
rect 201 478 203 480
rect 211 499 213 501
rect 211 492 213 494
rect 227 485 229 487
rect 227 478 229 480
rect 247 493 249 495
rect 258 493 260 495
rect 294 499 296 501
rect 278 485 280 487
rect 278 478 280 480
rect 294 492 296 494
rect 322 492 324 494
rect 332 492 334 494
rect 332 485 334 487
rect 342 490 344 492
rect 304 478 306 480
rect 362 492 364 494
rect 381 499 383 501
rect 410 478 412 480
rect 420 499 422 501
rect 420 492 422 494
rect 436 485 438 487
rect 436 478 438 480
rect 476 499 478 501
rect 456 493 458 495
rect 493 489 495 491
rect 510 499 512 501
rect 466 477 468 479
rect 540 499 542 501
rect 557 489 559 491
rect 574 499 576 501
rect 530 477 532 479
rect 604 499 606 501
rect 621 489 623 491
rect 638 499 640 501
rect 594 477 596 479
rect 9 379 11 381
rect 29 394 31 396
rect 29 387 31 389
rect 45 380 47 382
rect 45 373 47 375
rect 55 394 57 396
rect 73 380 75 382
rect 83 387 85 389
rect 83 380 85 382
rect 93 382 95 384
rect 113 379 115 381
rect 133 394 135 396
rect 133 387 135 389
rect 149 380 151 382
rect 149 373 151 375
rect 159 394 161 396
rect 177 380 179 382
rect 187 387 189 389
rect 187 380 189 382
rect 197 382 199 384
rect 217 380 219 382
rect 258 379 260 381
rect 236 373 238 375
rect 278 394 280 396
rect 278 387 280 389
rect 294 380 296 382
rect 294 373 296 375
rect 304 394 306 396
rect 322 380 324 382
rect 332 387 334 389
rect 332 380 334 382
rect 342 382 344 384
rect 362 380 364 382
rect 410 394 412 396
rect 381 373 383 375
rect 420 380 422 382
rect 436 394 438 396
rect 436 387 438 389
rect 420 373 422 375
rect 466 395 468 397
rect 530 395 532 397
rect 456 379 458 381
rect 476 373 478 375
rect 493 383 495 385
rect 510 373 512 375
rect 594 395 596 397
rect 540 373 542 375
rect 557 383 559 385
rect 574 373 576 375
rect 604 373 606 375
rect 621 383 623 385
rect 638 373 640 375
rect 20 355 22 357
rect 39 348 41 350
rect 59 346 61 348
rect 69 348 71 350
rect 69 341 71 343
rect 79 348 81 350
rect 97 334 99 336
rect 107 355 109 357
rect 107 348 109 350
rect 123 341 125 343
rect 123 334 125 336
rect 143 349 145 351
rect 163 346 165 348
rect 173 348 175 350
rect 173 341 175 343
rect 183 348 185 350
rect 201 334 203 336
rect 211 355 213 357
rect 211 348 213 350
rect 227 341 229 343
rect 227 334 229 336
rect 247 349 249 351
rect 258 349 260 351
rect 294 355 296 357
rect 278 341 280 343
rect 278 334 280 336
rect 294 348 296 350
rect 322 348 324 350
rect 332 348 334 350
rect 332 341 334 343
rect 342 346 344 348
rect 304 334 306 336
rect 362 348 364 350
rect 381 355 383 357
rect 410 334 412 336
rect 420 355 422 357
rect 420 348 422 350
rect 436 341 438 343
rect 436 334 438 336
rect 476 355 478 357
rect 456 349 458 351
rect 493 345 495 347
rect 510 355 512 357
rect 466 333 468 335
rect 540 355 542 357
rect 557 345 559 347
rect 574 355 576 357
rect 530 333 532 335
rect 604 355 606 357
rect 621 345 623 347
rect 638 355 640 357
rect 594 333 596 335
rect 9 235 11 237
rect 29 250 31 252
rect 29 243 31 245
rect 45 236 47 238
rect 45 229 47 231
rect 55 250 57 252
rect 73 236 75 238
rect 83 243 85 245
rect 83 236 85 238
rect 93 238 95 240
rect 113 235 115 237
rect 133 250 135 252
rect 133 243 135 245
rect 149 236 151 238
rect 149 229 151 231
rect 159 250 161 252
rect 177 236 179 238
rect 187 243 189 245
rect 187 236 189 238
rect 197 238 199 240
rect 217 236 219 238
rect 258 235 260 237
rect 236 229 238 231
rect 278 250 280 252
rect 278 243 280 245
rect 294 236 296 238
rect 294 229 296 231
rect 304 250 306 252
rect 322 236 324 238
rect 332 243 334 245
rect 332 236 334 238
rect 342 238 344 240
rect 362 236 364 238
rect 410 250 412 252
rect 381 229 383 231
rect 420 236 422 238
rect 436 250 438 252
rect 436 243 438 245
rect 420 229 422 231
rect 466 251 468 253
rect 530 251 532 253
rect 456 235 458 237
rect 476 229 478 231
rect 493 239 495 241
rect 510 229 512 231
rect 594 251 596 253
rect 540 229 542 231
rect 557 239 559 241
rect 574 229 576 231
rect 604 229 606 231
rect 621 239 623 241
rect 638 229 640 231
rect 20 211 22 213
rect 39 204 41 206
rect 59 202 61 204
rect 69 204 71 206
rect 69 197 71 199
rect 79 204 81 206
rect 97 190 99 192
rect 107 211 109 213
rect 107 204 109 206
rect 123 197 125 199
rect 123 190 125 192
rect 143 205 145 207
rect 163 202 165 204
rect 173 204 175 206
rect 173 197 175 199
rect 183 204 185 206
rect 201 190 203 192
rect 211 211 213 213
rect 211 204 213 206
rect 227 197 229 199
rect 227 190 229 192
rect 247 205 249 207
rect 258 205 260 207
rect 294 211 296 213
rect 278 197 280 199
rect 278 190 280 192
rect 294 204 296 206
rect 322 204 324 206
rect 332 204 334 206
rect 332 197 334 199
rect 342 202 344 204
rect 304 190 306 192
rect 362 204 364 206
rect 381 211 383 213
rect 410 190 412 192
rect 420 211 422 213
rect 420 204 422 206
rect 436 197 438 199
rect 436 190 438 192
rect 476 211 478 213
rect 456 205 458 207
rect 493 201 495 203
rect 510 211 512 213
rect 466 189 468 191
rect 540 211 542 213
rect 557 201 559 203
rect 574 211 576 213
rect 530 189 532 191
rect 604 211 606 213
rect 621 201 623 203
rect 638 211 640 213
rect 594 189 596 191
rect 9 91 11 93
rect 29 106 31 108
rect 29 99 31 101
rect 45 92 47 94
rect 45 85 47 87
rect 55 106 57 108
rect 73 92 75 94
rect 83 99 85 101
rect 83 92 85 94
rect 93 94 95 96
rect 113 91 115 93
rect 133 106 135 108
rect 133 99 135 101
rect 149 92 151 94
rect 149 85 151 87
rect 159 106 161 108
rect 177 92 179 94
rect 187 99 189 101
rect 187 92 189 94
rect 197 94 199 96
rect 217 92 219 94
rect 258 91 260 93
rect 236 85 238 87
rect 278 106 280 108
rect 278 99 280 101
rect 294 92 296 94
rect 294 85 296 87
rect 304 106 306 108
rect 322 92 324 94
rect 332 99 334 101
rect 332 92 334 94
rect 342 94 344 96
rect 362 92 364 94
rect 410 106 412 108
rect 381 85 383 87
rect 420 92 422 94
rect 436 106 438 108
rect 436 99 438 101
rect 420 85 422 87
rect 466 107 468 109
rect 530 107 532 109
rect 456 91 458 93
rect 476 85 478 87
rect 493 95 495 97
rect 510 85 512 87
rect 594 107 596 109
rect 540 85 542 87
rect 557 95 559 97
rect 574 85 576 87
rect 604 85 606 87
rect 621 95 623 97
rect 638 85 640 87
rect 20 67 22 69
rect 39 60 41 62
rect 59 58 61 60
rect 69 60 71 62
rect 69 53 71 55
rect 79 60 81 62
rect 97 46 99 48
rect 107 67 109 69
rect 107 60 109 62
rect 123 53 125 55
rect 123 46 125 48
rect 143 61 145 63
rect 163 58 165 60
rect 173 60 175 62
rect 173 53 175 55
rect 183 60 185 62
rect 201 46 203 48
rect 211 67 213 69
rect 211 60 213 62
rect 227 53 229 55
rect 227 46 229 48
rect 247 61 249 63
rect 258 61 260 63
rect 294 67 296 69
rect 278 53 280 55
rect 278 46 280 48
rect 294 60 296 62
rect 322 60 324 62
rect 332 60 334 62
rect 332 53 334 55
rect 342 58 344 60
rect 304 46 306 48
rect 362 60 364 62
rect 381 67 383 69
rect 410 46 412 48
rect 420 67 422 69
rect 420 60 422 62
rect 436 53 438 55
rect 436 46 438 48
rect 476 67 478 69
rect 456 61 458 63
rect 493 57 495 59
rect 510 67 512 69
rect 466 45 468 47
rect 540 67 542 69
rect 557 57 559 59
rect 574 67 576 69
rect 530 45 532 47
rect 604 67 606 69
rect 621 57 623 59
rect 638 67 640 69
rect 594 45 596 47
<< pdifct1 >>
rect 19 531 21 533
rect 103 538 105 540
rect 103 531 105 533
rect 123 531 125 533
rect 207 538 209 540
rect 207 531 209 533
rect 247 534 249 536
rect 247 527 249 529
rect 268 531 270 533
rect 352 538 354 540
rect 352 531 354 533
rect 392 534 394 536
rect 392 527 394 529
rect 446 531 448 533
rect 520 524 522 526
rect 584 524 586 526
rect 648 524 650 526
rect 9 489 11 491
rect 9 482 11 484
rect 49 485 51 487
rect 49 478 51 480
rect 133 485 135 487
rect 153 485 155 487
rect 153 478 155 480
rect 237 485 239 487
rect 268 485 270 487
rect 352 485 354 487
rect 352 478 354 480
rect 392 489 394 491
rect 392 482 394 484
rect 446 485 448 487
rect 520 492 522 494
rect 584 492 586 494
rect 648 492 650 494
rect 19 387 21 389
rect 103 394 105 396
rect 103 387 105 389
rect 123 387 125 389
rect 207 394 209 396
rect 207 387 209 389
rect 247 390 249 392
rect 247 383 249 385
rect 268 387 270 389
rect 352 394 354 396
rect 352 387 354 389
rect 392 390 394 392
rect 392 383 394 385
rect 446 387 448 389
rect 520 380 522 382
rect 584 380 586 382
rect 648 380 650 382
rect 9 345 11 347
rect 9 338 11 340
rect 49 341 51 343
rect 49 334 51 336
rect 133 341 135 343
rect 153 341 155 343
rect 153 334 155 336
rect 237 341 239 343
rect 268 341 270 343
rect 352 341 354 343
rect 352 334 354 336
rect 392 345 394 347
rect 392 338 394 340
rect 446 341 448 343
rect 520 348 522 350
rect 584 348 586 350
rect 648 348 650 350
rect 19 243 21 245
rect 103 250 105 252
rect 103 243 105 245
rect 123 243 125 245
rect 207 250 209 252
rect 207 243 209 245
rect 247 246 249 248
rect 247 239 249 241
rect 268 243 270 245
rect 352 250 354 252
rect 352 243 354 245
rect 392 246 394 248
rect 392 239 394 241
rect 446 243 448 245
rect 520 236 522 238
rect 584 236 586 238
rect 648 236 650 238
rect 9 201 11 203
rect 9 194 11 196
rect 49 197 51 199
rect 49 190 51 192
rect 133 197 135 199
rect 153 197 155 199
rect 153 190 155 192
rect 237 197 239 199
rect 268 197 270 199
rect 352 197 354 199
rect 352 190 354 192
rect 392 201 394 203
rect 392 194 394 196
rect 446 197 448 199
rect 520 204 522 206
rect 584 204 586 206
rect 648 204 650 206
rect 19 99 21 101
rect 103 106 105 108
rect 103 99 105 101
rect 123 99 125 101
rect 207 106 209 108
rect 207 99 209 101
rect 247 102 249 104
rect 247 95 249 97
rect 268 99 270 101
rect 352 106 354 108
rect 352 99 354 101
rect 392 102 394 104
rect 392 95 394 97
rect 446 99 448 101
rect 520 92 522 94
rect 584 92 586 94
rect 648 92 650 94
rect 9 57 11 59
rect 9 50 11 52
rect 49 53 51 55
rect 49 46 51 48
rect 133 53 135 55
rect 153 53 155 55
rect 153 46 155 48
rect 237 53 239 55
rect 268 53 270 55
rect 352 53 354 55
rect 352 46 354 48
rect 392 57 394 59
rect 392 50 394 52
rect 446 53 448 55
rect 520 60 522 62
rect 584 60 586 62
rect 648 60 650 62
<< alu0 >>
rect 47 567 53 573
rect 36 564 40 566
rect 47 565 49 567
rect 51 565 53 567
rect 47 564 53 565
rect 71 566 91 567
rect 71 564 73 566
rect 75 564 91 566
rect 36 562 37 564
rect 39 562 40 564
rect 71 563 91 564
rect 36 559 40 562
rect 16 555 40 559
rect 16 551 20 555
rect 62 559 66 561
rect 62 557 63 559
rect 65 557 66 559
rect 15 549 20 551
rect 15 547 16 549
rect 18 547 20 549
rect 24 550 40 551
rect 24 548 26 550
rect 28 548 40 550
rect 24 547 40 548
rect 15 545 20 547
rect 16 543 20 545
rect 16 540 32 543
rect 16 539 29 540
rect 28 538 29 539
rect 31 538 32 540
rect 28 533 32 538
rect 28 531 29 533
rect 31 531 32 533
rect 28 529 32 531
rect 36 541 40 547
rect 62 551 66 557
rect 55 547 66 551
rect 87 559 91 563
rect 151 567 157 573
rect 215 572 221 573
rect 215 570 217 572
rect 219 570 221 572
rect 215 569 221 570
rect 234 572 240 573
rect 234 570 236 572
rect 238 570 240 572
rect 234 569 240 570
rect 102 560 103 562
rect 87 555 99 559
rect 95 550 99 555
rect 95 548 96 550
rect 98 548 99 550
rect 55 541 59 547
rect 36 540 59 541
rect 36 538 55 540
rect 57 538 59 540
rect 36 537 59 538
rect 36 526 40 537
rect 95 536 99 548
rect 82 533 99 536
rect 82 531 83 533
rect 85 532 99 533
rect 85 531 86 532
rect 7 525 40 526
rect 7 523 9 525
rect 11 523 40 525
rect 7 522 40 523
rect 44 526 48 528
rect 44 524 45 526
rect 47 524 48 526
rect 44 519 48 524
rect 71 526 77 527
rect 71 524 73 526
rect 75 524 77 526
rect 44 517 45 519
rect 47 517 48 519
rect 71 517 77 524
rect 82 526 86 531
rect 140 564 144 566
rect 151 565 153 567
rect 155 565 157 567
rect 151 564 157 565
rect 175 566 195 567
rect 175 564 177 566
rect 179 564 195 566
rect 140 562 141 564
rect 143 562 144 564
rect 175 563 195 564
rect 140 559 144 562
rect 120 555 144 559
rect 120 551 124 555
rect 166 559 170 561
rect 166 557 167 559
rect 169 557 170 559
rect 119 549 124 551
rect 119 547 120 549
rect 122 547 124 549
rect 128 550 144 551
rect 128 548 130 550
rect 132 548 144 550
rect 128 547 144 548
rect 119 545 124 547
rect 120 543 124 545
rect 120 540 136 543
rect 120 539 133 540
rect 132 538 133 539
rect 135 538 136 540
rect 132 533 136 538
rect 132 531 133 533
rect 135 531 136 533
rect 132 529 136 531
rect 140 541 144 547
rect 166 551 170 557
rect 159 547 170 551
rect 191 559 195 563
rect 296 567 302 573
rect 360 572 366 573
rect 360 570 362 572
rect 364 570 366 572
rect 360 569 366 570
rect 379 572 385 573
rect 379 570 381 572
rect 383 570 385 572
rect 379 569 385 570
rect 206 560 207 562
rect 191 555 203 559
rect 199 550 203 555
rect 199 548 200 550
rect 202 548 203 550
rect 159 541 163 547
rect 140 540 163 541
rect 140 538 159 540
rect 161 538 163 540
rect 140 537 163 538
rect 82 524 83 526
rect 85 524 86 526
rect 82 522 86 524
rect 91 528 97 529
rect 91 526 93 528
rect 95 526 97 528
rect 140 526 144 537
rect 199 536 203 548
rect 285 564 289 566
rect 296 565 298 567
rect 300 565 302 567
rect 296 564 302 565
rect 320 566 340 567
rect 320 564 322 566
rect 324 564 340 566
rect 225 559 243 560
rect 225 557 227 559
rect 229 557 243 559
rect 225 556 243 557
rect 239 550 243 556
rect 239 548 240 550
rect 242 548 243 550
rect 218 543 224 544
rect 186 533 203 536
rect 186 531 187 533
rect 189 532 203 533
rect 189 531 190 532
rect 91 517 97 526
rect 111 525 144 526
rect 111 523 113 525
rect 115 523 144 525
rect 111 522 144 523
rect 148 526 152 528
rect 148 524 149 526
rect 151 524 152 526
rect 148 519 152 524
rect 175 526 181 527
rect 175 524 177 526
rect 179 524 181 526
rect 148 517 149 519
rect 151 517 152 519
rect 175 517 181 524
rect 186 526 190 531
rect 239 535 243 548
rect 228 531 243 535
rect 186 524 187 526
rect 189 524 190 526
rect 186 522 190 524
rect 195 528 201 529
rect 195 526 197 528
rect 199 526 201 528
rect 228 527 232 531
rect 246 527 247 538
rect 285 562 286 564
rect 288 562 289 564
rect 320 563 340 564
rect 285 559 289 562
rect 265 555 289 559
rect 265 551 269 555
rect 311 559 315 561
rect 311 557 312 559
rect 314 557 315 559
rect 264 549 269 551
rect 264 547 265 549
rect 267 547 269 549
rect 273 550 289 551
rect 273 548 275 550
rect 277 548 289 550
rect 273 547 289 548
rect 264 545 269 547
rect 265 543 269 545
rect 265 540 281 543
rect 265 539 278 540
rect 277 538 278 539
rect 280 538 281 540
rect 277 533 281 538
rect 277 531 278 533
rect 280 531 281 533
rect 277 529 281 531
rect 285 541 289 547
rect 311 551 315 557
rect 304 547 315 551
rect 336 559 340 563
rect 414 567 420 573
rect 414 565 416 567
rect 418 565 420 567
rect 414 564 420 565
rect 427 564 431 566
rect 351 560 352 562
rect 336 555 348 559
rect 344 550 348 555
rect 344 548 345 550
rect 347 548 348 550
rect 304 541 308 547
rect 285 540 308 541
rect 285 538 304 540
rect 306 538 308 540
rect 285 537 308 538
rect 195 517 201 526
rect 215 526 232 527
rect 215 524 217 526
rect 219 524 232 526
rect 215 523 232 524
rect 285 526 289 537
rect 344 536 348 548
rect 427 562 428 564
rect 430 562 431 564
rect 370 559 388 560
rect 370 557 372 559
rect 374 557 388 559
rect 370 556 388 557
rect 384 550 388 556
rect 384 548 385 550
rect 387 548 388 550
rect 363 543 369 544
rect 331 533 348 536
rect 331 531 332 533
rect 334 532 348 533
rect 334 531 335 532
rect 256 525 289 526
rect 256 523 258 525
rect 260 523 289 525
rect 256 522 289 523
rect 293 526 297 528
rect 293 524 294 526
rect 296 524 297 526
rect 234 519 240 520
rect 234 517 236 519
rect 238 517 240 519
rect 293 519 297 524
rect 320 526 326 527
rect 320 524 322 526
rect 324 524 326 526
rect 293 517 294 519
rect 296 517 297 519
rect 320 517 326 524
rect 331 526 335 531
rect 384 535 388 548
rect 401 559 405 561
rect 401 557 402 559
rect 404 557 405 559
rect 401 551 405 557
rect 427 559 431 562
rect 427 555 451 559
rect 401 547 412 551
rect 373 531 388 535
rect 331 524 332 526
rect 334 524 335 526
rect 331 522 335 524
rect 340 528 346 529
rect 340 526 342 528
rect 344 526 346 528
rect 373 527 377 531
rect 391 527 392 538
rect 340 517 346 526
rect 360 526 377 527
rect 360 524 362 526
rect 364 524 377 526
rect 360 523 377 524
rect 408 541 412 547
rect 447 551 451 555
rect 427 550 443 551
rect 427 548 439 550
rect 441 548 443 550
rect 427 547 443 548
rect 447 549 452 551
rect 447 547 449 549
rect 451 547 452 549
rect 427 541 431 547
rect 447 545 452 547
rect 447 543 451 545
rect 408 540 431 541
rect 408 538 410 540
rect 412 538 431 540
rect 408 537 431 538
rect 419 526 423 528
rect 419 524 420 526
rect 422 524 423 526
rect 379 519 385 520
rect 379 517 381 519
rect 383 517 385 519
rect 419 519 423 524
rect 427 526 431 537
rect 435 540 451 543
rect 435 538 436 540
rect 438 539 451 540
rect 438 538 439 539
rect 435 533 439 538
rect 464 565 470 566
rect 464 563 466 565
rect 468 563 470 565
rect 464 562 470 563
rect 474 565 480 573
rect 474 563 476 565
rect 478 563 480 565
rect 491 567 506 568
rect 491 565 493 567
rect 495 565 506 567
rect 491 564 506 565
rect 474 562 480 563
rect 464 542 468 562
rect 502 559 506 564
rect 509 567 513 573
rect 509 565 510 567
rect 512 565 513 567
rect 509 563 513 565
rect 488 556 499 558
rect 488 554 496 556
rect 498 554 499 556
rect 502 557 516 559
rect 502 555 517 557
rect 488 552 499 554
rect 512 553 514 555
rect 516 553 517 555
rect 488 542 492 552
rect 512 551 517 553
rect 464 541 492 542
rect 464 539 466 541
rect 468 540 492 541
rect 468 539 489 540
rect 464 538 489 539
rect 491 538 492 540
rect 508 541 509 547
rect 488 536 492 538
rect 435 531 436 533
rect 438 531 439 533
rect 435 529 439 531
rect 512 534 516 551
rect 500 530 516 534
rect 528 565 534 566
rect 528 563 530 565
rect 532 563 534 565
rect 528 562 534 563
rect 538 565 544 573
rect 538 563 540 565
rect 542 563 544 565
rect 555 567 570 568
rect 555 565 557 567
rect 559 565 570 567
rect 555 564 570 565
rect 538 562 544 563
rect 528 542 532 562
rect 566 559 570 564
rect 573 567 577 573
rect 573 565 574 567
rect 576 565 577 567
rect 573 563 577 565
rect 552 556 563 558
rect 552 554 560 556
rect 562 554 563 556
rect 566 557 580 559
rect 566 555 581 557
rect 552 552 563 554
rect 576 553 578 555
rect 580 553 581 555
rect 552 542 556 552
rect 576 551 581 553
rect 528 541 556 542
rect 528 539 530 541
rect 532 540 556 541
rect 532 539 553 540
rect 528 538 553 539
rect 555 538 556 540
rect 572 541 573 547
rect 552 536 556 538
rect 427 525 460 526
rect 427 523 456 525
rect 458 523 460 525
rect 427 522 460 523
rect 491 529 504 530
rect 491 527 493 529
rect 495 527 504 529
rect 491 526 504 527
rect 576 534 580 551
rect 564 530 580 534
rect 555 529 568 530
rect 555 527 557 529
rect 559 527 568 529
rect 592 565 598 566
rect 592 563 594 565
rect 596 563 598 565
rect 592 562 598 563
rect 602 565 608 573
rect 602 563 604 565
rect 606 563 608 565
rect 619 567 634 568
rect 619 565 621 567
rect 623 565 634 567
rect 619 564 634 565
rect 602 562 608 563
rect 592 542 596 562
rect 630 559 634 564
rect 637 567 641 573
rect 637 565 638 567
rect 640 565 641 567
rect 637 563 641 565
rect 616 556 627 558
rect 616 554 624 556
rect 626 554 627 556
rect 630 557 644 559
rect 630 555 645 557
rect 616 552 627 554
rect 640 553 642 555
rect 644 553 645 555
rect 616 542 620 552
rect 640 551 645 553
rect 592 541 620 542
rect 592 539 594 541
rect 596 540 620 541
rect 596 539 617 540
rect 592 538 617 539
rect 619 538 620 540
rect 636 541 637 547
rect 616 536 620 538
rect 555 526 568 527
rect 640 534 644 551
rect 628 530 644 534
rect 619 529 632 530
rect 619 527 621 529
rect 623 527 632 529
rect 619 526 632 527
rect 419 517 420 519
rect 422 517 423 519
rect 475 519 479 521
rect 475 517 476 519
rect 478 517 479 519
rect 508 519 514 520
rect 508 517 510 519
rect 512 517 514 519
rect 539 519 543 521
rect 539 517 540 519
rect 542 517 543 519
rect 572 519 578 520
rect 572 517 574 519
rect 576 517 578 519
rect 603 519 607 521
rect 603 517 604 519
rect 606 517 607 519
rect 636 519 642 520
rect 636 517 638 519
rect 640 517 642 519
rect 18 499 20 501
rect 22 499 24 501
rect 18 498 24 499
rect 26 494 43 495
rect 26 492 39 494
rect 41 492 43 494
rect 26 491 43 492
rect 57 492 63 501
rect 11 480 12 491
rect 26 487 30 491
rect 57 490 59 492
rect 61 490 63 492
rect 57 489 63 490
rect 68 494 72 496
rect 68 492 69 494
rect 71 492 72 494
rect 15 483 30 487
rect 15 470 19 483
rect 68 487 72 492
rect 77 494 83 501
rect 106 499 107 501
rect 109 499 110 501
rect 77 492 79 494
rect 81 492 83 494
rect 77 491 83 492
rect 106 494 110 499
rect 106 492 107 494
rect 109 492 110 494
rect 106 490 110 492
rect 114 495 147 496
rect 114 493 143 495
rect 145 493 147 495
rect 114 492 147 493
rect 161 492 167 501
rect 68 486 69 487
rect 55 485 69 486
rect 71 485 72 487
rect 55 482 72 485
rect 34 474 40 475
rect 15 468 16 470
rect 18 468 19 470
rect 15 462 19 468
rect 15 461 33 462
rect 15 459 29 461
rect 31 459 33 461
rect 15 458 33 459
rect 55 470 59 482
rect 114 481 118 492
rect 161 490 163 492
rect 165 490 167 492
rect 161 489 167 490
rect 172 494 176 496
rect 172 492 173 494
rect 175 492 176 494
rect 95 480 118 481
rect 95 478 97 480
rect 99 478 118 480
rect 95 477 118 478
rect 95 471 99 477
rect 55 468 56 470
rect 58 468 59 470
rect 55 463 59 468
rect 55 459 67 463
rect 51 456 52 458
rect 63 455 67 459
rect 88 467 99 471
rect 88 461 92 467
rect 114 471 118 477
rect 122 487 126 489
rect 122 485 123 487
rect 125 485 126 487
rect 122 480 126 485
rect 122 478 123 480
rect 125 479 126 480
rect 125 478 138 479
rect 122 475 138 478
rect 134 473 138 475
rect 134 471 139 473
rect 114 470 130 471
rect 114 468 126 470
rect 128 468 130 470
rect 114 467 130 468
rect 134 469 136 471
rect 138 469 139 471
rect 134 467 139 469
rect 88 459 89 461
rect 91 459 92 461
rect 88 457 92 459
rect 134 463 138 467
rect 114 459 138 463
rect 114 456 118 459
rect 63 454 83 455
rect 114 454 115 456
rect 117 454 118 456
rect 63 452 79 454
rect 81 452 83 454
rect 63 451 83 452
rect 101 453 107 454
rect 101 451 103 453
rect 105 451 107 453
rect 114 452 118 454
rect 172 487 176 492
rect 181 494 187 501
rect 210 499 211 501
rect 213 499 214 501
rect 181 492 183 494
rect 185 492 187 494
rect 181 491 187 492
rect 210 494 214 499
rect 293 499 294 501
rect 296 499 297 501
rect 210 492 211 494
rect 213 492 214 494
rect 210 490 214 492
rect 218 495 251 496
rect 218 493 247 495
rect 249 493 251 495
rect 218 492 251 493
rect 256 495 289 496
rect 256 493 258 495
rect 260 493 289 495
rect 256 492 289 493
rect 172 486 173 487
rect 159 485 173 486
rect 175 485 176 487
rect 159 482 176 485
rect 159 470 163 482
rect 218 481 222 492
rect 199 480 222 481
rect 199 478 201 480
rect 203 478 222 480
rect 199 477 222 478
rect 199 471 203 477
rect 159 468 160 470
rect 162 468 163 470
rect 159 463 163 468
rect 159 459 171 463
rect 155 456 156 458
rect 18 448 24 449
rect 18 446 20 448
rect 22 446 24 448
rect 18 445 24 446
rect 37 448 43 449
rect 37 446 39 448
rect 41 446 43 448
rect 37 445 43 446
rect 101 445 107 451
rect 167 455 171 459
rect 192 467 203 471
rect 192 461 196 467
rect 218 471 222 477
rect 226 487 230 489
rect 226 485 227 487
rect 229 485 230 487
rect 226 480 230 485
rect 226 478 227 480
rect 229 479 230 480
rect 229 478 242 479
rect 226 475 242 478
rect 238 473 242 475
rect 238 471 243 473
rect 218 470 234 471
rect 218 468 230 470
rect 232 468 234 470
rect 218 467 234 468
rect 238 469 240 471
rect 242 469 243 471
rect 238 467 243 469
rect 192 459 193 461
rect 195 459 196 461
rect 192 457 196 459
rect 238 463 242 467
rect 218 459 242 463
rect 218 456 222 459
rect 167 454 187 455
rect 218 454 219 456
rect 221 454 222 456
rect 167 452 183 454
rect 185 452 187 454
rect 167 451 187 452
rect 205 453 211 454
rect 205 451 207 453
rect 209 451 211 453
rect 218 452 222 454
rect 277 487 281 489
rect 277 485 278 487
rect 280 485 281 487
rect 277 480 281 485
rect 277 479 278 480
rect 265 478 278 479
rect 280 478 281 480
rect 265 475 281 478
rect 285 481 289 492
rect 293 494 297 499
rect 293 492 294 494
rect 296 492 297 494
rect 293 490 297 492
rect 320 494 326 501
rect 320 492 322 494
rect 324 492 326 494
rect 320 491 326 492
rect 331 494 335 496
rect 331 492 332 494
rect 334 492 335 494
rect 285 480 308 481
rect 285 478 304 480
rect 306 478 308 480
rect 285 477 308 478
rect 265 473 269 475
rect 264 471 269 473
rect 285 471 289 477
rect 264 469 265 471
rect 267 469 269 471
rect 264 467 269 469
rect 273 470 289 471
rect 273 468 275 470
rect 277 468 289 470
rect 273 467 289 468
rect 265 463 269 467
rect 304 471 308 477
rect 331 487 335 492
rect 340 492 346 501
rect 379 499 381 501
rect 383 499 385 501
rect 379 498 385 499
rect 419 499 420 501
rect 422 499 423 501
rect 340 490 342 492
rect 344 490 346 492
rect 360 494 377 495
rect 360 492 362 494
rect 364 492 377 494
rect 360 491 377 492
rect 340 489 346 490
rect 331 485 332 487
rect 334 486 335 487
rect 334 485 348 486
rect 331 482 348 485
rect 304 467 315 471
rect 265 459 289 463
rect 285 456 289 459
rect 311 461 315 467
rect 311 459 312 461
rect 314 459 315 461
rect 311 457 315 459
rect 344 470 348 482
rect 344 468 345 470
rect 347 468 348 470
rect 344 463 348 468
rect 336 459 348 463
rect 285 454 286 456
rect 288 454 289 456
rect 336 455 340 459
rect 351 456 352 458
rect 373 487 377 491
rect 373 483 388 487
rect 363 474 369 475
rect 384 470 388 483
rect 391 480 392 491
rect 384 468 385 470
rect 387 468 388 470
rect 384 462 388 468
rect 419 494 423 499
rect 475 499 476 501
rect 478 499 479 501
rect 475 497 479 499
rect 508 499 510 501
rect 512 499 514 501
rect 508 498 514 499
rect 539 499 540 501
rect 542 499 543 501
rect 539 497 543 499
rect 572 499 574 501
rect 576 499 578 501
rect 572 498 578 499
rect 603 499 604 501
rect 606 499 607 501
rect 603 497 607 499
rect 636 499 638 501
rect 640 499 642 501
rect 636 498 642 499
rect 419 492 420 494
rect 422 492 423 494
rect 419 490 423 492
rect 427 495 460 496
rect 427 493 456 495
rect 458 493 460 495
rect 427 492 460 493
rect 427 481 431 492
rect 408 480 431 481
rect 408 478 410 480
rect 412 478 431 480
rect 408 477 431 478
rect 408 471 412 477
rect 370 461 388 462
rect 370 459 372 461
rect 374 459 388 461
rect 370 458 388 459
rect 401 467 412 471
rect 401 461 405 467
rect 427 471 431 477
rect 435 487 439 489
rect 491 491 504 492
rect 491 489 493 491
rect 495 489 504 491
rect 491 488 504 489
rect 435 485 436 487
rect 438 485 439 487
rect 435 480 439 485
rect 500 484 516 488
rect 435 478 436 480
rect 438 479 439 480
rect 438 478 451 479
rect 435 475 451 478
rect 447 473 451 475
rect 447 471 452 473
rect 427 470 443 471
rect 427 468 439 470
rect 441 468 443 470
rect 427 467 443 468
rect 447 469 449 471
rect 451 469 452 471
rect 447 467 452 469
rect 401 459 402 461
rect 404 459 405 461
rect 401 457 405 459
rect 447 463 451 467
rect 427 459 451 463
rect 488 480 492 482
rect 320 454 340 455
rect 285 452 289 454
rect 296 453 302 454
rect 296 451 298 453
rect 300 451 302 453
rect 320 452 322 454
rect 324 452 340 454
rect 320 451 340 452
rect 427 456 431 459
rect 427 454 428 456
rect 430 454 431 456
rect 205 445 211 451
rect 296 445 302 451
rect 414 453 420 454
rect 414 451 416 453
rect 418 451 420 453
rect 427 452 431 454
rect 464 479 489 480
rect 464 477 466 479
rect 468 478 489 479
rect 491 478 492 480
rect 468 477 492 478
rect 464 476 492 477
rect 464 456 468 476
rect 488 466 492 476
rect 508 471 509 477
rect 512 467 516 484
rect 488 464 499 466
rect 488 462 496 464
rect 498 462 499 464
rect 512 465 517 467
rect 512 463 514 465
rect 516 463 517 465
rect 488 460 499 462
rect 502 461 517 463
rect 502 459 516 461
rect 464 455 470 456
rect 464 453 466 455
rect 468 453 470 455
rect 464 452 470 453
rect 474 455 480 456
rect 474 453 476 455
rect 478 453 480 455
rect 502 454 506 459
rect 555 491 568 492
rect 555 489 557 491
rect 559 489 568 491
rect 555 488 568 489
rect 564 484 580 488
rect 552 480 556 482
rect 360 448 366 449
rect 360 446 362 448
rect 364 446 366 448
rect 360 445 366 446
rect 379 448 385 449
rect 379 446 381 448
rect 383 446 385 448
rect 379 445 385 446
rect 414 445 420 451
rect 474 445 480 453
rect 491 453 506 454
rect 491 451 493 453
rect 495 451 506 453
rect 491 450 506 451
rect 509 453 513 455
rect 509 451 510 453
rect 512 451 513 453
rect 528 479 553 480
rect 528 477 530 479
rect 532 478 553 479
rect 555 478 556 480
rect 532 477 556 478
rect 528 476 556 477
rect 528 456 532 476
rect 552 466 556 476
rect 572 471 573 477
rect 576 467 580 484
rect 552 464 563 466
rect 552 462 560 464
rect 562 462 563 464
rect 576 465 581 467
rect 576 463 578 465
rect 580 463 581 465
rect 552 460 563 462
rect 566 461 581 463
rect 619 491 632 492
rect 619 489 621 491
rect 623 489 632 491
rect 619 488 632 489
rect 628 484 644 488
rect 616 480 620 482
rect 566 459 580 461
rect 528 455 534 456
rect 528 453 530 455
rect 532 453 534 455
rect 528 452 534 453
rect 538 455 544 456
rect 538 453 540 455
rect 542 453 544 455
rect 566 454 570 459
rect 509 445 513 451
rect 538 445 544 453
rect 555 453 570 454
rect 555 451 557 453
rect 559 451 570 453
rect 555 450 570 451
rect 573 453 577 455
rect 573 451 574 453
rect 576 451 577 453
rect 592 479 617 480
rect 592 477 594 479
rect 596 478 617 479
rect 619 478 620 480
rect 596 477 620 478
rect 592 476 620 477
rect 592 456 596 476
rect 616 466 620 476
rect 636 471 637 477
rect 640 467 644 484
rect 616 464 627 466
rect 616 462 624 464
rect 626 462 627 464
rect 640 465 645 467
rect 640 463 642 465
rect 644 463 645 465
rect 616 460 627 462
rect 630 461 645 463
rect 630 459 644 461
rect 592 455 598 456
rect 592 453 594 455
rect 596 453 598 455
rect 592 452 598 453
rect 602 455 608 456
rect 602 453 604 455
rect 606 453 608 455
rect 630 454 634 459
rect 573 445 577 451
rect 602 445 608 453
rect 619 453 634 454
rect 619 451 621 453
rect 623 451 634 453
rect 619 450 634 451
rect 637 453 641 455
rect 637 451 638 453
rect 640 451 641 453
rect 637 445 641 451
rect 47 423 53 429
rect 36 420 40 422
rect 47 421 49 423
rect 51 421 53 423
rect 47 420 53 421
rect 71 422 91 423
rect 71 420 73 422
rect 75 420 91 422
rect 36 418 37 420
rect 39 418 40 420
rect 71 419 91 420
rect 36 415 40 418
rect 16 411 40 415
rect 16 407 20 411
rect 62 415 66 417
rect 62 413 63 415
rect 65 413 66 415
rect 15 405 20 407
rect 15 403 16 405
rect 18 403 20 405
rect 24 406 40 407
rect 24 404 26 406
rect 28 404 40 406
rect 24 403 40 404
rect 15 401 20 403
rect 16 399 20 401
rect 16 396 32 399
rect 16 395 29 396
rect 28 394 29 395
rect 31 394 32 396
rect 28 389 32 394
rect 28 387 29 389
rect 31 387 32 389
rect 28 385 32 387
rect 36 397 40 403
rect 62 407 66 413
rect 55 403 66 407
rect 87 415 91 419
rect 151 423 157 429
rect 215 428 221 429
rect 215 426 217 428
rect 219 426 221 428
rect 215 425 221 426
rect 234 428 240 429
rect 234 426 236 428
rect 238 426 240 428
rect 234 425 240 426
rect 102 416 103 418
rect 87 411 99 415
rect 95 406 99 411
rect 95 404 96 406
rect 98 404 99 406
rect 55 397 59 403
rect 36 396 59 397
rect 36 394 55 396
rect 57 394 59 396
rect 36 393 59 394
rect 36 382 40 393
rect 95 392 99 404
rect 82 389 99 392
rect 82 387 83 389
rect 85 388 99 389
rect 85 387 86 388
rect 7 381 40 382
rect 7 379 9 381
rect 11 379 40 381
rect 7 378 40 379
rect 44 382 48 384
rect 44 380 45 382
rect 47 380 48 382
rect 44 375 48 380
rect 71 382 77 383
rect 71 380 73 382
rect 75 380 77 382
rect 44 373 45 375
rect 47 373 48 375
rect 71 373 77 380
rect 82 382 86 387
rect 140 420 144 422
rect 151 421 153 423
rect 155 421 157 423
rect 151 420 157 421
rect 175 422 195 423
rect 175 420 177 422
rect 179 420 195 422
rect 140 418 141 420
rect 143 418 144 420
rect 175 419 195 420
rect 140 415 144 418
rect 120 411 144 415
rect 120 407 124 411
rect 166 415 170 417
rect 166 413 167 415
rect 169 413 170 415
rect 119 405 124 407
rect 119 403 120 405
rect 122 403 124 405
rect 128 406 144 407
rect 128 404 130 406
rect 132 404 144 406
rect 128 403 144 404
rect 119 401 124 403
rect 120 399 124 401
rect 120 396 136 399
rect 120 395 133 396
rect 132 394 133 395
rect 135 394 136 396
rect 132 389 136 394
rect 132 387 133 389
rect 135 387 136 389
rect 132 385 136 387
rect 140 397 144 403
rect 166 407 170 413
rect 159 403 170 407
rect 191 415 195 419
rect 296 423 302 429
rect 360 428 366 429
rect 360 426 362 428
rect 364 426 366 428
rect 360 425 366 426
rect 379 428 385 429
rect 379 426 381 428
rect 383 426 385 428
rect 379 425 385 426
rect 206 416 207 418
rect 191 411 203 415
rect 199 406 203 411
rect 199 404 200 406
rect 202 404 203 406
rect 159 397 163 403
rect 140 396 163 397
rect 140 394 159 396
rect 161 394 163 396
rect 140 393 163 394
rect 82 380 83 382
rect 85 380 86 382
rect 82 378 86 380
rect 91 384 97 385
rect 91 382 93 384
rect 95 382 97 384
rect 140 382 144 393
rect 199 392 203 404
rect 285 420 289 422
rect 296 421 298 423
rect 300 421 302 423
rect 296 420 302 421
rect 320 422 340 423
rect 320 420 322 422
rect 324 420 340 422
rect 225 415 243 416
rect 225 413 227 415
rect 229 413 243 415
rect 225 412 243 413
rect 239 406 243 412
rect 239 404 240 406
rect 242 404 243 406
rect 218 399 224 400
rect 186 389 203 392
rect 186 387 187 389
rect 189 388 203 389
rect 189 387 190 388
rect 91 373 97 382
rect 111 381 144 382
rect 111 379 113 381
rect 115 379 144 381
rect 111 378 144 379
rect 148 382 152 384
rect 148 380 149 382
rect 151 380 152 382
rect 148 375 152 380
rect 175 382 181 383
rect 175 380 177 382
rect 179 380 181 382
rect 148 373 149 375
rect 151 373 152 375
rect 175 373 181 380
rect 186 382 190 387
rect 239 391 243 404
rect 228 387 243 391
rect 186 380 187 382
rect 189 380 190 382
rect 186 378 190 380
rect 195 384 201 385
rect 195 382 197 384
rect 199 382 201 384
rect 228 383 232 387
rect 246 383 247 394
rect 285 418 286 420
rect 288 418 289 420
rect 320 419 340 420
rect 285 415 289 418
rect 265 411 289 415
rect 265 407 269 411
rect 311 415 315 417
rect 311 413 312 415
rect 314 413 315 415
rect 264 405 269 407
rect 264 403 265 405
rect 267 403 269 405
rect 273 406 289 407
rect 273 404 275 406
rect 277 404 289 406
rect 273 403 289 404
rect 264 401 269 403
rect 265 399 269 401
rect 265 396 281 399
rect 265 395 278 396
rect 277 394 278 395
rect 280 394 281 396
rect 277 389 281 394
rect 277 387 278 389
rect 280 387 281 389
rect 277 385 281 387
rect 285 397 289 403
rect 311 407 315 413
rect 304 403 315 407
rect 336 415 340 419
rect 414 423 420 429
rect 414 421 416 423
rect 418 421 420 423
rect 414 420 420 421
rect 427 420 431 422
rect 351 416 352 418
rect 336 411 348 415
rect 344 406 348 411
rect 344 404 345 406
rect 347 404 348 406
rect 304 397 308 403
rect 285 396 308 397
rect 285 394 304 396
rect 306 394 308 396
rect 285 393 308 394
rect 195 373 201 382
rect 215 382 232 383
rect 215 380 217 382
rect 219 380 232 382
rect 215 379 232 380
rect 285 382 289 393
rect 344 392 348 404
rect 427 418 428 420
rect 430 418 431 420
rect 370 415 388 416
rect 370 413 372 415
rect 374 413 388 415
rect 370 412 388 413
rect 384 406 388 412
rect 384 404 385 406
rect 387 404 388 406
rect 363 399 369 400
rect 331 389 348 392
rect 331 387 332 389
rect 334 388 348 389
rect 334 387 335 388
rect 256 381 289 382
rect 256 379 258 381
rect 260 379 289 381
rect 256 378 289 379
rect 293 382 297 384
rect 293 380 294 382
rect 296 380 297 382
rect 234 375 240 376
rect 234 373 236 375
rect 238 373 240 375
rect 293 375 297 380
rect 320 382 326 383
rect 320 380 322 382
rect 324 380 326 382
rect 293 373 294 375
rect 296 373 297 375
rect 320 373 326 380
rect 331 382 335 387
rect 384 391 388 404
rect 401 415 405 417
rect 401 413 402 415
rect 404 413 405 415
rect 401 407 405 413
rect 427 415 431 418
rect 427 411 451 415
rect 401 403 412 407
rect 373 387 388 391
rect 331 380 332 382
rect 334 380 335 382
rect 331 378 335 380
rect 340 384 346 385
rect 340 382 342 384
rect 344 382 346 384
rect 373 383 377 387
rect 391 383 392 394
rect 340 373 346 382
rect 360 382 377 383
rect 360 380 362 382
rect 364 380 377 382
rect 360 379 377 380
rect 408 397 412 403
rect 447 407 451 411
rect 427 406 443 407
rect 427 404 439 406
rect 441 404 443 406
rect 427 403 443 404
rect 447 405 452 407
rect 447 403 449 405
rect 451 403 452 405
rect 427 397 431 403
rect 447 401 452 403
rect 447 399 451 401
rect 408 396 431 397
rect 408 394 410 396
rect 412 394 431 396
rect 408 393 431 394
rect 419 382 423 384
rect 419 380 420 382
rect 422 380 423 382
rect 379 375 385 376
rect 379 373 381 375
rect 383 373 385 375
rect 419 375 423 380
rect 427 382 431 393
rect 435 396 451 399
rect 435 394 436 396
rect 438 395 451 396
rect 438 394 439 395
rect 435 389 439 394
rect 464 421 470 422
rect 464 419 466 421
rect 468 419 470 421
rect 464 418 470 419
rect 474 421 480 429
rect 474 419 476 421
rect 478 419 480 421
rect 491 423 506 424
rect 491 421 493 423
rect 495 421 506 423
rect 491 420 506 421
rect 474 418 480 419
rect 464 398 468 418
rect 502 415 506 420
rect 509 423 513 429
rect 509 421 510 423
rect 512 421 513 423
rect 509 419 513 421
rect 488 412 499 414
rect 488 410 496 412
rect 498 410 499 412
rect 502 413 516 415
rect 502 411 517 413
rect 488 408 499 410
rect 512 409 514 411
rect 516 409 517 411
rect 488 398 492 408
rect 512 407 517 409
rect 464 397 492 398
rect 464 395 466 397
rect 468 396 492 397
rect 468 395 489 396
rect 464 394 489 395
rect 491 394 492 396
rect 508 397 509 403
rect 488 392 492 394
rect 435 387 436 389
rect 438 387 439 389
rect 435 385 439 387
rect 512 390 516 407
rect 500 386 516 390
rect 528 421 534 422
rect 528 419 530 421
rect 532 419 534 421
rect 528 418 534 419
rect 538 421 544 429
rect 538 419 540 421
rect 542 419 544 421
rect 555 423 570 424
rect 555 421 557 423
rect 559 421 570 423
rect 555 420 570 421
rect 538 418 544 419
rect 528 398 532 418
rect 566 415 570 420
rect 573 423 577 429
rect 573 421 574 423
rect 576 421 577 423
rect 573 419 577 421
rect 552 412 563 414
rect 552 410 560 412
rect 562 410 563 412
rect 566 413 580 415
rect 566 411 581 413
rect 552 408 563 410
rect 576 409 578 411
rect 580 409 581 411
rect 552 398 556 408
rect 576 407 581 409
rect 528 397 556 398
rect 528 395 530 397
rect 532 396 556 397
rect 532 395 553 396
rect 528 394 553 395
rect 555 394 556 396
rect 572 397 573 403
rect 552 392 556 394
rect 427 381 460 382
rect 427 379 456 381
rect 458 379 460 381
rect 427 378 460 379
rect 491 385 504 386
rect 491 383 493 385
rect 495 383 504 385
rect 491 382 504 383
rect 576 390 580 407
rect 564 386 580 390
rect 555 385 568 386
rect 555 383 557 385
rect 559 383 568 385
rect 592 421 598 422
rect 592 419 594 421
rect 596 419 598 421
rect 592 418 598 419
rect 602 421 608 429
rect 602 419 604 421
rect 606 419 608 421
rect 619 423 634 424
rect 619 421 621 423
rect 623 421 634 423
rect 619 420 634 421
rect 602 418 608 419
rect 592 398 596 418
rect 630 415 634 420
rect 637 423 641 429
rect 637 421 638 423
rect 640 421 641 423
rect 637 419 641 421
rect 616 412 627 414
rect 616 410 624 412
rect 626 410 627 412
rect 630 413 644 415
rect 630 411 645 413
rect 616 408 627 410
rect 640 409 642 411
rect 644 409 645 411
rect 616 398 620 408
rect 640 407 645 409
rect 592 397 620 398
rect 592 395 594 397
rect 596 396 620 397
rect 596 395 617 396
rect 592 394 617 395
rect 619 394 620 396
rect 636 397 637 403
rect 616 392 620 394
rect 555 382 568 383
rect 640 390 644 407
rect 628 386 644 390
rect 619 385 632 386
rect 619 383 621 385
rect 623 383 632 385
rect 619 382 632 383
rect 419 373 420 375
rect 422 373 423 375
rect 475 375 479 377
rect 475 373 476 375
rect 478 373 479 375
rect 508 375 514 376
rect 508 373 510 375
rect 512 373 514 375
rect 539 375 543 377
rect 539 373 540 375
rect 542 373 543 375
rect 572 375 578 376
rect 572 373 574 375
rect 576 373 578 375
rect 603 375 607 377
rect 603 373 604 375
rect 606 373 607 375
rect 636 375 642 376
rect 636 373 638 375
rect 640 373 642 375
rect 18 355 20 357
rect 22 355 24 357
rect 18 354 24 355
rect 26 350 43 351
rect 26 348 39 350
rect 41 348 43 350
rect 26 347 43 348
rect 57 348 63 357
rect 11 336 12 347
rect 26 343 30 347
rect 57 346 59 348
rect 61 346 63 348
rect 57 345 63 346
rect 68 350 72 352
rect 68 348 69 350
rect 71 348 72 350
rect 15 339 30 343
rect 15 326 19 339
rect 68 343 72 348
rect 77 350 83 357
rect 106 355 107 357
rect 109 355 110 357
rect 77 348 79 350
rect 81 348 83 350
rect 77 347 83 348
rect 106 350 110 355
rect 106 348 107 350
rect 109 348 110 350
rect 106 346 110 348
rect 114 351 147 352
rect 114 349 143 351
rect 145 349 147 351
rect 114 348 147 349
rect 161 348 167 357
rect 68 342 69 343
rect 55 341 69 342
rect 71 341 72 343
rect 55 338 72 341
rect 34 330 40 331
rect 15 324 16 326
rect 18 324 19 326
rect 15 318 19 324
rect 15 317 33 318
rect 15 315 29 317
rect 31 315 33 317
rect 15 314 33 315
rect 55 326 59 338
rect 114 337 118 348
rect 161 346 163 348
rect 165 346 167 348
rect 161 345 167 346
rect 172 350 176 352
rect 172 348 173 350
rect 175 348 176 350
rect 95 336 118 337
rect 95 334 97 336
rect 99 334 118 336
rect 95 333 118 334
rect 95 327 99 333
rect 55 324 56 326
rect 58 324 59 326
rect 55 319 59 324
rect 55 315 67 319
rect 51 312 52 314
rect 63 311 67 315
rect 88 323 99 327
rect 88 317 92 323
rect 114 327 118 333
rect 122 343 126 345
rect 122 341 123 343
rect 125 341 126 343
rect 122 336 126 341
rect 122 334 123 336
rect 125 335 126 336
rect 125 334 138 335
rect 122 331 138 334
rect 134 329 138 331
rect 134 327 139 329
rect 114 326 130 327
rect 114 324 126 326
rect 128 324 130 326
rect 114 323 130 324
rect 134 325 136 327
rect 138 325 139 327
rect 134 323 139 325
rect 88 315 89 317
rect 91 315 92 317
rect 88 313 92 315
rect 134 319 138 323
rect 114 315 138 319
rect 114 312 118 315
rect 63 310 83 311
rect 114 310 115 312
rect 117 310 118 312
rect 63 308 79 310
rect 81 308 83 310
rect 63 307 83 308
rect 101 309 107 310
rect 101 307 103 309
rect 105 307 107 309
rect 114 308 118 310
rect 172 343 176 348
rect 181 350 187 357
rect 210 355 211 357
rect 213 355 214 357
rect 181 348 183 350
rect 185 348 187 350
rect 181 347 187 348
rect 210 350 214 355
rect 293 355 294 357
rect 296 355 297 357
rect 210 348 211 350
rect 213 348 214 350
rect 210 346 214 348
rect 218 351 251 352
rect 218 349 247 351
rect 249 349 251 351
rect 218 348 251 349
rect 256 351 289 352
rect 256 349 258 351
rect 260 349 289 351
rect 256 348 289 349
rect 172 342 173 343
rect 159 341 173 342
rect 175 341 176 343
rect 159 338 176 341
rect 159 326 163 338
rect 218 337 222 348
rect 199 336 222 337
rect 199 334 201 336
rect 203 334 222 336
rect 199 333 222 334
rect 199 327 203 333
rect 159 324 160 326
rect 162 324 163 326
rect 159 319 163 324
rect 159 315 171 319
rect 155 312 156 314
rect 18 304 24 305
rect 18 302 20 304
rect 22 302 24 304
rect 18 301 24 302
rect 37 304 43 305
rect 37 302 39 304
rect 41 302 43 304
rect 37 301 43 302
rect 101 301 107 307
rect 167 311 171 315
rect 192 323 203 327
rect 192 317 196 323
rect 218 327 222 333
rect 226 343 230 345
rect 226 341 227 343
rect 229 341 230 343
rect 226 336 230 341
rect 226 334 227 336
rect 229 335 230 336
rect 229 334 242 335
rect 226 331 242 334
rect 238 329 242 331
rect 238 327 243 329
rect 218 326 234 327
rect 218 324 230 326
rect 232 324 234 326
rect 218 323 234 324
rect 238 325 240 327
rect 242 325 243 327
rect 238 323 243 325
rect 192 315 193 317
rect 195 315 196 317
rect 192 313 196 315
rect 238 319 242 323
rect 218 315 242 319
rect 218 312 222 315
rect 167 310 187 311
rect 218 310 219 312
rect 221 310 222 312
rect 167 308 183 310
rect 185 308 187 310
rect 167 307 187 308
rect 205 309 211 310
rect 205 307 207 309
rect 209 307 211 309
rect 218 308 222 310
rect 277 343 281 345
rect 277 341 278 343
rect 280 341 281 343
rect 277 336 281 341
rect 277 335 278 336
rect 265 334 278 335
rect 280 334 281 336
rect 265 331 281 334
rect 285 337 289 348
rect 293 350 297 355
rect 293 348 294 350
rect 296 348 297 350
rect 293 346 297 348
rect 320 350 326 357
rect 320 348 322 350
rect 324 348 326 350
rect 320 347 326 348
rect 331 350 335 352
rect 331 348 332 350
rect 334 348 335 350
rect 285 336 308 337
rect 285 334 304 336
rect 306 334 308 336
rect 285 333 308 334
rect 265 329 269 331
rect 264 327 269 329
rect 285 327 289 333
rect 264 325 265 327
rect 267 325 269 327
rect 264 323 269 325
rect 273 326 289 327
rect 273 324 275 326
rect 277 324 289 326
rect 273 323 289 324
rect 265 319 269 323
rect 304 327 308 333
rect 331 343 335 348
rect 340 348 346 357
rect 379 355 381 357
rect 383 355 385 357
rect 379 354 385 355
rect 419 355 420 357
rect 422 355 423 357
rect 340 346 342 348
rect 344 346 346 348
rect 360 350 377 351
rect 360 348 362 350
rect 364 348 377 350
rect 360 347 377 348
rect 340 345 346 346
rect 331 341 332 343
rect 334 342 335 343
rect 334 341 348 342
rect 331 338 348 341
rect 304 323 315 327
rect 265 315 289 319
rect 285 312 289 315
rect 311 317 315 323
rect 311 315 312 317
rect 314 315 315 317
rect 311 313 315 315
rect 344 326 348 338
rect 344 324 345 326
rect 347 324 348 326
rect 344 319 348 324
rect 336 315 348 319
rect 285 310 286 312
rect 288 310 289 312
rect 336 311 340 315
rect 351 312 352 314
rect 373 343 377 347
rect 373 339 388 343
rect 363 330 369 331
rect 384 326 388 339
rect 391 336 392 347
rect 384 324 385 326
rect 387 324 388 326
rect 384 318 388 324
rect 419 350 423 355
rect 475 355 476 357
rect 478 355 479 357
rect 475 353 479 355
rect 508 355 510 357
rect 512 355 514 357
rect 508 354 514 355
rect 539 355 540 357
rect 542 355 543 357
rect 539 353 543 355
rect 572 355 574 357
rect 576 355 578 357
rect 572 354 578 355
rect 603 355 604 357
rect 606 355 607 357
rect 603 353 607 355
rect 636 355 638 357
rect 640 355 642 357
rect 636 354 642 355
rect 419 348 420 350
rect 422 348 423 350
rect 419 346 423 348
rect 427 351 460 352
rect 427 349 456 351
rect 458 349 460 351
rect 427 348 460 349
rect 427 337 431 348
rect 408 336 431 337
rect 408 334 410 336
rect 412 334 431 336
rect 408 333 431 334
rect 408 327 412 333
rect 370 317 388 318
rect 370 315 372 317
rect 374 315 388 317
rect 370 314 388 315
rect 401 323 412 327
rect 401 317 405 323
rect 427 327 431 333
rect 435 343 439 345
rect 491 347 504 348
rect 491 345 493 347
rect 495 345 504 347
rect 491 344 504 345
rect 435 341 436 343
rect 438 341 439 343
rect 435 336 439 341
rect 500 340 516 344
rect 435 334 436 336
rect 438 335 439 336
rect 438 334 451 335
rect 435 331 451 334
rect 447 329 451 331
rect 447 327 452 329
rect 427 326 443 327
rect 427 324 439 326
rect 441 324 443 326
rect 427 323 443 324
rect 447 325 449 327
rect 451 325 452 327
rect 447 323 452 325
rect 401 315 402 317
rect 404 315 405 317
rect 401 313 405 315
rect 447 319 451 323
rect 427 315 451 319
rect 488 336 492 338
rect 320 310 340 311
rect 285 308 289 310
rect 296 309 302 310
rect 296 307 298 309
rect 300 307 302 309
rect 320 308 322 310
rect 324 308 340 310
rect 320 307 340 308
rect 427 312 431 315
rect 427 310 428 312
rect 430 310 431 312
rect 205 301 211 307
rect 296 301 302 307
rect 414 309 420 310
rect 414 307 416 309
rect 418 307 420 309
rect 427 308 431 310
rect 464 335 489 336
rect 464 333 466 335
rect 468 334 489 335
rect 491 334 492 336
rect 468 333 492 334
rect 464 332 492 333
rect 464 312 468 332
rect 488 322 492 332
rect 508 327 509 333
rect 512 323 516 340
rect 488 320 499 322
rect 488 318 496 320
rect 498 318 499 320
rect 512 321 517 323
rect 512 319 514 321
rect 516 319 517 321
rect 488 316 499 318
rect 502 317 517 319
rect 502 315 516 317
rect 464 311 470 312
rect 464 309 466 311
rect 468 309 470 311
rect 464 308 470 309
rect 474 311 480 312
rect 474 309 476 311
rect 478 309 480 311
rect 502 310 506 315
rect 555 347 568 348
rect 555 345 557 347
rect 559 345 568 347
rect 555 344 568 345
rect 564 340 580 344
rect 552 336 556 338
rect 360 304 366 305
rect 360 302 362 304
rect 364 302 366 304
rect 360 301 366 302
rect 379 304 385 305
rect 379 302 381 304
rect 383 302 385 304
rect 379 301 385 302
rect 414 301 420 307
rect 474 301 480 309
rect 491 309 506 310
rect 491 307 493 309
rect 495 307 506 309
rect 491 306 506 307
rect 509 309 513 311
rect 509 307 510 309
rect 512 307 513 309
rect 528 335 553 336
rect 528 333 530 335
rect 532 334 553 335
rect 555 334 556 336
rect 532 333 556 334
rect 528 332 556 333
rect 528 312 532 332
rect 552 322 556 332
rect 572 327 573 333
rect 576 323 580 340
rect 552 320 563 322
rect 552 318 560 320
rect 562 318 563 320
rect 576 321 581 323
rect 576 319 578 321
rect 580 319 581 321
rect 552 316 563 318
rect 566 317 581 319
rect 619 347 632 348
rect 619 345 621 347
rect 623 345 632 347
rect 619 344 632 345
rect 628 340 644 344
rect 616 336 620 338
rect 566 315 580 317
rect 528 311 534 312
rect 528 309 530 311
rect 532 309 534 311
rect 528 308 534 309
rect 538 311 544 312
rect 538 309 540 311
rect 542 309 544 311
rect 566 310 570 315
rect 509 301 513 307
rect 538 301 544 309
rect 555 309 570 310
rect 555 307 557 309
rect 559 307 570 309
rect 555 306 570 307
rect 573 309 577 311
rect 573 307 574 309
rect 576 307 577 309
rect 592 335 617 336
rect 592 333 594 335
rect 596 334 617 335
rect 619 334 620 336
rect 596 333 620 334
rect 592 332 620 333
rect 592 312 596 332
rect 616 322 620 332
rect 636 327 637 333
rect 640 323 644 340
rect 616 320 627 322
rect 616 318 624 320
rect 626 318 627 320
rect 640 321 645 323
rect 640 319 642 321
rect 644 319 645 321
rect 616 316 627 318
rect 630 317 645 319
rect 630 315 644 317
rect 592 311 598 312
rect 592 309 594 311
rect 596 309 598 311
rect 592 308 598 309
rect 602 311 608 312
rect 602 309 604 311
rect 606 309 608 311
rect 630 310 634 315
rect 573 301 577 307
rect 602 301 608 309
rect 619 309 634 310
rect 619 307 621 309
rect 623 307 634 309
rect 619 306 634 307
rect 637 309 641 311
rect 637 307 638 309
rect 640 307 641 309
rect 637 301 641 307
rect 47 279 53 285
rect 36 276 40 278
rect 47 277 49 279
rect 51 277 53 279
rect 47 276 53 277
rect 71 278 91 279
rect 71 276 73 278
rect 75 276 91 278
rect 36 274 37 276
rect 39 274 40 276
rect 71 275 91 276
rect 36 271 40 274
rect 16 267 40 271
rect 16 263 20 267
rect 62 271 66 273
rect 62 269 63 271
rect 65 269 66 271
rect 15 261 20 263
rect 15 259 16 261
rect 18 259 20 261
rect 24 262 40 263
rect 24 260 26 262
rect 28 260 40 262
rect 24 259 40 260
rect 15 257 20 259
rect 16 255 20 257
rect 16 252 32 255
rect 16 251 29 252
rect 28 250 29 251
rect 31 250 32 252
rect 28 245 32 250
rect 28 243 29 245
rect 31 243 32 245
rect 28 241 32 243
rect 36 253 40 259
rect 62 263 66 269
rect 55 259 66 263
rect 87 271 91 275
rect 151 279 157 285
rect 215 284 221 285
rect 215 282 217 284
rect 219 282 221 284
rect 215 281 221 282
rect 234 284 240 285
rect 234 282 236 284
rect 238 282 240 284
rect 234 281 240 282
rect 102 272 103 274
rect 87 267 99 271
rect 95 262 99 267
rect 95 260 96 262
rect 98 260 99 262
rect 55 253 59 259
rect 36 252 59 253
rect 36 250 55 252
rect 57 250 59 252
rect 36 249 59 250
rect 36 238 40 249
rect 95 248 99 260
rect 82 245 99 248
rect 82 243 83 245
rect 85 244 99 245
rect 85 243 86 244
rect 7 237 40 238
rect 7 235 9 237
rect 11 235 40 237
rect 7 234 40 235
rect 44 238 48 240
rect 44 236 45 238
rect 47 236 48 238
rect 44 231 48 236
rect 71 238 77 239
rect 71 236 73 238
rect 75 236 77 238
rect 44 229 45 231
rect 47 229 48 231
rect 71 229 77 236
rect 82 238 86 243
rect 140 276 144 278
rect 151 277 153 279
rect 155 277 157 279
rect 151 276 157 277
rect 175 278 195 279
rect 175 276 177 278
rect 179 276 195 278
rect 140 274 141 276
rect 143 274 144 276
rect 175 275 195 276
rect 140 271 144 274
rect 120 267 144 271
rect 120 263 124 267
rect 166 271 170 273
rect 166 269 167 271
rect 169 269 170 271
rect 119 261 124 263
rect 119 259 120 261
rect 122 259 124 261
rect 128 262 144 263
rect 128 260 130 262
rect 132 260 144 262
rect 128 259 144 260
rect 119 257 124 259
rect 120 255 124 257
rect 120 252 136 255
rect 120 251 133 252
rect 132 250 133 251
rect 135 250 136 252
rect 132 245 136 250
rect 132 243 133 245
rect 135 243 136 245
rect 132 241 136 243
rect 140 253 144 259
rect 166 263 170 269
rect 159 259 170 263
rect 191 271 195 275
rect 296 279 302 285
rect 360 284 366 285
rect 360 282 362 284
rect 364 282 366 284
rect 360 281 366 282
rect 379 284 385 285
rect 379 282 381 284
rect 383 282 385 284
rect 379 281 385 282
rect 206 272 207 274
rect 191 267 203 271
rect 199 262 203 267
rect 199 260 200 262
rect 202 260 203 262
rect 159 253 163 259
rect 140 252 163 253
rect 140 250 159 252
rect 161 250 163 252
rect 140 249 163 250
rect 82 236 83 238
rect 85 236 86 238
rect 82 234 86 236
rect 91 240 97 241
rect 91 238 93 240
rect 95 238 97 240
rect 140 238 144 249
rect 199 248 203 260
rect 285 276 289 278
rect 296 277 298 279
rect 300 277 302 279
rect 296 276 302 277
rect 320 278 340 279
rect 320 276 322 278
rect 324 276 340 278
rect 225 271 243 272
rect 225 269 227 271
rect 229 269 243 271
rect 225 268 243 269
rect 239 262 243 268
rect 239 260 240 262
rect 242 260 243 262
rect 218 255 224 256
rect 186 245 203 248
rect 186 243 187 245
rect 189 244 203 245
rect 189 243 190 244
rect 91 229 97 238
rect 111 237 144 238
rect 111 235 113 237
rect 115 235 144 237
rect 111 234 144 235
rect 148 238 152 240
rect 148 236 149 238
rect 151 236 152 238
rect 148 231 152 236
rect 175 238 181 239
rect 175 236 177 238
rect 179 236 181 238
rect 148 229 149 231
rect 151 229 152 231
rect 175 229 181 236
rect 186 238 190 243
rect 239 247 243 260
rect 228 243 243 247
rect 186 236 187 238
rect 189 236 190 238
rect 186 234 190 236
rect 195 240 201 241
rect 195 238 197 240
rect 199 238 201 240
rect 228 239 232 243
rect 246 239 247 250
rect 285 274 286 276
rect 288 274 289 276
rect 320 275 340 276
rect 285 271 289 274
rect 265 267 289 271
rect 265 263 269 267
rect 311 271 315 273
rect 311 269 312 271
rect 314 269 315 271
rect 264 261 269 263
rect 264 259 265 261
rect 267 259 269 261
rect 273 262 289 263
rect 273 260 275 262
rect 277 260 289 262
rect 273 259 289 260
rect 264 257 269 259
rect 265 255 269 257
rect 265 252 281 255
rect 265 251 278 252
rect 277 250 278 251
rect 280 250 281 252
rect 277 245 281 250
rect 277 243 278 245
rect 280 243 281 245
rect 277 241 281 243
rect 285 253 289 259
rect 311 263 315 269
rect 304 259 315 263
rect 336 271 340 275
rect 414 279 420 285
rect 414 277 416 279
rect 418 277 420 279
rect 414 276 420 277
rect 427 276 431 278
rect 351 272 352 274
rect 336 267 348 271
rect 344 262 348 267
rect 344 260 345 262
rect 347 260 348 262
rect 304 253 308 259
rect 285 252 308 253
rect 285 250 304 252
rect 306 250 308 252
rect 285 249 308 250
rect 195 229 201 238
rect 215 238 232 239
rect 215 236 217 238
rect 219 236 232 238
rect 215 235 232 236
rect 285 238 289 249
rect 344 248 348 260
rect 427 274 428 276
rect 430 274 431 276
rect 370 271 388 272
rect 370 269 372 271
rect 374 269 388 271
rect 370 268 388 269
rect 384 262 388 268
rect 384 260 385 262
rect 387 260 388 262
rect 363 255 369 256
rect 331 245 348 248
rect 331 243 332 245
rect 334 244 348 245
rect 334 243 335 244
rect 256 237 289 238
rect 256 235 258 237
rect 260 235 289 237
rect 256 234 289 235
rect 293 238 297 240
rect 293 236 294 238
rect 296 236 297 238
rect 234 231 240 232
rect 234 229 236 231
rect 238 229 240 231
rect 293 231 297 236
rect 320 238 326 239
rect 320 236 322 238
rect 324 236 326 238
rect 293 229 294 231
rect 296 229 297 231
rect 320 229 326 236
rect 331 238 335 243
rect 384 247 388 260
rect 401 271 405 273
rect 401 269 402 271
rect 404 269 405 271
rect 401 263 405 269
rect 427 271 431 274
rect 427 267 451 271
rect 401 259 412 263
rect 373 243 388 247
rect 331 236 332 238
rect 334 236 335 238
rect 331 234 335 236
rect 340 240 346 241
rect 340 238 342 240
rect 344 238 346 240
rect 373 239 377 243
rect 391 239 392 250
rect 340 229 346 238
rect 360 238 377 239
rect 360 236 362 238
rect 364 236 377 238
rect 360 235 377 236
rect 408 253 412 259
rect 447 263 451 267
rect 427 262 443 263
rect 427 260 439 262
rect 441 260 443 262
rect 427 259 443 260
rect 447 261 452 263
rect 447 259 449 261
rect 451 259 452 261
rect 427 253 431 259
rect 447 257 452 259
rect 447 255 451 257
rect 408 252 431 253
rect 408 250 410 252
rect 412 250 431 252
rect 408 249 431 250
rect 419 238 423 240
rect 419 236 420 238
rect 422 236 423 238
rect 379 231 385 232
rect 379 229 381 231
rect 383 229 385 231
rect 419 231 423 236
rect 427 238 431 249
rect 435 252 451 255
rect 435 250 436 252
rect 438 251 451 252
rect 438 250 439 251
rect 435 245 439 250
rect 464 277 470 278
rect 464 275 466 277
rect 468 275 470 277
rect 464 274 470 275
rect 474 277 480 285
rect 474 275 476 277
rect 478 275 480 277
rect 491 279 506 280
rect 491 277 493 279
rect 495 277 506 279
rect 491 276 506 277
rect 474 274 480 275
rect 464 254 468 274
rect 502 271 506 276
rect 509 279 513 285
rect 509 277 510 279
rect 512 277 513 279
rect 509 275 513 277
rect 488 268 499 270
rect 488 266 496 268
rect 498 266 499 268
rect 502 269 516 271
rect 502 267 517 269
rect 488 264 499 266
rect 512 265 514 267
rect 516 265 517 267
rect 488 254 492 264
rect 512 263 517 265
rect 464 253 492 254
rect 464 251 466 253
rect 468 252 492 253
rect 468 251 489 252
rect 464 250 489 251
rect 491 250 492 252
rect 508 253 509 259
rect 488 248 492 250
rect 435 243 436 245
rect 438 243 439 245
rect 435 241 439 243
rect 512 246 516 263
rect 500 242 516 246
rect 528 277 534 278
rect 528 275 530 277
rect 532 275 534 277
rect 528 274 534 275
rect 538 277 544 285
rect 538 275 540 277
rect 542 275 544 277
rect 555 279 570 280
rect 555 277 557 279
rect 559 277 570 279
rect 555 276 570 277
rect 538 274 544 275
rect 528 254 532 274
rect 566 271 570 276
rect 573 279 577 285
rect 573 277 574 279
rect 576 277 577 279
rect 573 275 577 277
rect 552 268 563 270
rect 552 266 560 268
rect 562 266 563 268
rect 566 269 580 271
rect 566 267 581 269
rect 552 264 563 266
rect 576 265 578 267
rect 580 265 581 267
rect 552 254 556 264
rect 576 263 581 265
rect 528 253 556 254
rect 528 251 530 253
rect 532 252 556 253
rect 532 251 553 252
rect 528 250 553 251
rect 555 250 556 252
rect 572 253 573 259
rect 552 248 556 250
rect 427 237 460 238
rect 427 235 456 237
rect 458 235 460 237
rect 427 234 460 235
rect 491 241 504 242
rect 491 239 493 241
rect 495 239 504 241
rect 491 238 504 239
rect 576 246 580 263
rect 564 242 580 246
rect 555 241 568 242
rect 555 239 557 241
rect 559 239 568 241
rect 592 277 598 278
rect 592 275 594 277
rect 596 275 598 277
rect 592 274 598 275
rect 602 277 608 285
rect 602 275 604 277
rect 606 275 608 277
rect 619 279 634 280
rect 619 277 621 279
rect 623 277 634 279
rect 619 276 634 277
rect 602 274 608 275
rect 592 254 596 274
rect 630 271 634 276
rect 637 279 641 285
rect 637 277 638 279
rect 640 277 641 279
rect 637 275 641 277
rect 616 268 627 270
rect 616 266 624 268
rect 626 266 627 268
rect 630 269 644 271
rect 630 267 645 269
rect 616 264 627 266
rect 640 265 642 267
rect 644 265 645 267
rect 616 254 620 264
rect 640 263 645 265
rect 592 253 620 254
rect 592 251 594 253
rect 596 252 620 253
rect 596 251 617 252
rect 592 250 617 251
rect 619 250 620 252
rect 636 253 637 259
rect 616 248 620 250
rect 555 238 568 239
rect 640 246 644 263
rect 628 242 644 246
rect 619 241 632 242
rect 619 239 621 241
rect 623 239 632 241
rect 619 238 632 239
rect 419 229 420 231
rect 422 229 423 231
rect 475 231 479 233
rect 475 229 476 231
rect 478 229 479 231
rect 508 231 514 232
rect 508 229 510 231
rect 512 229 514 231
rect 539 231 543 233
rect 539 229 540 231
rect 542 229 543 231
rect 572 231 578 232
rect 572 229 574 231
rect 576 229 578 231
rect 603 231 607 233
rect 603 229 604 231
rect 606 229 607 231
rect 636 231 642 232
rect 636 229 638 231
rect 640 229 642 231
rect 18 211 20 213
rect 22 211 24 213
rect 18 210 24 211
rect 26 206 43 207
rect 26 204 39 206
rect 41 204 43 206
rect 26 203 43 204
rect 57 204 63 213
rect 11 192 12 203
rect 26 199 30 203
rect 57 202 59 204
rect 61 202 63 204
rect 57 201 63 202
rect 68 206 72 208
rect 68 204 69 206
rect 71 204 72 206
rect 15 195 30 199
rect 15 182 19 195
rect 68 199 72 204
rect 77 206 83 213
rect 106 211 107 213
rect 109 211 110 213
rect 77 204 79 206
rect 81 204 83 206
rect 77 203 83 204
rect 106 206 110 211
rect 106 204 107 206
rect 109 204 110 206
rect 106 202 110 204
rect 114 207 147 208
rect 114 205 143 207
rect 145 205 147 207
rect 114 204 147 205
rect 161 204 167 213
rect 68 198 69 199
rect 55 197 69 198
rect 71 197 72 199
rect 55 194 72 197
rect 34 186 40 187
rect 15 180 16 182
rect 18 180 19 182
rect 15 174 19 180
rect 15 173 33 174
rect 15 171 29 173
rect 31 171 33 173
rect 15 170 33 171
rect 55 182 59 194
rect 114 193 118 204
rect 161 202 163 204
rect 165 202 167 204
rect 161 201 167 202
rect 172 206 176 208
rect 172 204 173 206
rect 175 204 176 206
rect 95 192 118 193
rect 95 190 97 192
rect 99 190 118 192
rect 95 189 118 190
rect 95 183 99 189
rect 55 180 56 182
rect 58 180 59 182
rect 55 175 59 180
rect 55 171 67 175
rect 51 168 52 170
rect 63 167 67 171
rect 88 179 99 183
rect 88 173 92 179
rect 114 183 118 189
rect 122 199 126 201
rect 122 197 123 199
rect 125 197 126 199
rect 122 192 126 197
rect 122 190 123 192
rect 125 191 126 192
rect 125 190 138 191
rect 122 187 138 190
rect 134 185 138 187
rect 134 183 139 185
rect 114 182 130 183
rect 114 180 126 182
rect 128 180 130 182
rect 114 179 130 180
rect 134 181 136 183
rect 138 181 139 183
rect 134 179 139 181
rect 88 171 89 173
rect 91 171 92 173
rect 88 169 92 171
rect 134 175 138 179
rect 114 171 138 175
rect 114 168 118 171
rect 63 166 83 167
rect 114 166 115 168
rect 117 166 118 168
rect 63 164 79 166
rect 81 164 83 166
rect 63 163 83 164
rect 101 165 107 166
rect 101 163 103 165
rect 105 163 107 165
rect 114 164 118 166
rect 172 199 176 204
rect 181 206 187 213
rect 210 211 211 213
rect 213 211 214 213
rect 181 204 183 206
rect 185 204 187 206
rect 181 203 187 204
rect 210 206 214 211
rect 293 211 294 213
rect 296 211 297 213
rect 210 204 211 206
rect 213 204 214 206
rect 210 202 214 204
rect 218 207 251 208
rect 218 205 247 207
rect 249 205 251 207
rect 218 204 251 205
rect 256 207 289 208
rect 256 205 258 207
rect 260 205 289 207
rect 256 204 289 205
rect 172 198 173 199
rect 159 197 173 198
rect 175 197 176 199
rect 159 194 176 197
rect 159 182 163 194
rect 218 193 222 204
rect 199 192 222 193
rect 199 190 201 192
rect 203 190 222 192
rect 199 189 222 190
rect 199 183 203 189
rect 159 180 160 182
rect 162 180 163 182
rect 159 175 163 180
rect 159 171 171 175
rect 155 168 156 170
rect 18 160 24 161
rect 18 158 20 160
rect 22 158 24 160
rect 18 157 24 158
rect 37 160 43 161
rect 37 158 39 160
rect 41 158 43 160
rect 37 157 43 158
rect 101 157 107 163
rect 167 167 171 171
rect 192 179 203 183
rect 192 173 196 179
rect 218 183 222 189
rect 226 199 230 201
rect 226 197 227 199
rect 229 197 230 199
rect 226 192 230 197
rect 226 190 227 192
rect 229 191 230 192
rect 229 190 242 191
rect 226 187 242 190
rect 238 185 242 187
rect 238 183 243 185
rect 218 182 234 183
rect 218 180 230 182
rect 232 180 234 182
rect 218 179 234 180
rect 238 181 240 183
rect 242 181 243 183
rect 238 179 243 181
rect 192 171 193 173
rect 195 171 196 173
rect 192 169 196 171
rect 238 175 242 179
rect 218 171 242 175
rect 218 168 222 171
rect 167 166 187 167
rect 218 166 219 168
rect 221 166 222 168
rect 167 164 183 166
rect 185 164 187 166
rect 167 163 187 164
rect 205 165 211 166
rect 205 163 207 165
rect 209 163 211 165
rect 218 164 222 166
rect 277 199 281 201
rect 277 197 278 199
rect 280 197 281 199
rect 277 192 281 197
rect 277 191 278 192
rect 265 190 278 191
rect 280 190 281 192
rect 265 187 281 190
rect 285 193 289 204
rect 293 206 297 211
rect 293 204 294 206
rect 296 204 297 206
rect 293 202 297 204
rect 320 206 326 213
rect 320 204 322 206
rect 324 204 326 206
rect 320 203 326 204
rect 331 206 335 208
rect 331 204 332 206
rect 334 204 335 206
rect 285 192 308 193
rect 285 190 304 192
rect 306 190 308 192
rect 285 189 308 190
rect 265 185 269 187
rect 264 183 269 185
rect 285 183 289 189
rect 264 181 265 183
rect 267 181 269 183
rect 264 179 269 181
rect 273 182 289 183
rect 273 180 275 182
rect 277 180 289 182
rect 273 179 289 180
rect 265 175 269 179
rect 304 183 308 189
rect 331 199 335 204
rect 340 204 346 213
rect 379 211 381 213
rect 383 211 385 213
rect 379 210 385 211
rect 419 211 420 213
rect 422 211 423 213
rect 340 202 342 204
rect 344 202 346 204
rect 360 206 377 207
rect 360 204 362 206
rect 364 204 377 206
rect 360 203 377 204
rect 340 201 346 202
rect 331 197 332 199
rect 334 198 335 199
rect 334 197 348 198
rect 331 194 348 197
rect 304 179 315 183
rect 265 171 289 175
rect 285 168 289 171
rect 311 173 315 179
rect 311 171 312 173
rect 314 171 315 173
rect 311 169 315 171
rect 344 182 348 194
rect 344 180 345 182
rect 347 180 348 182
rect 344 175 348 180
rect 336 171 348 175
rect 285 166 286 168
rect 288 166 289 168
rect 336 167 340 171
rect 351 168 352 170
rect 373 199 377 203
rect 373 195 388 199
rect 363 186 369 187
rect 384 182 388 195
rect 391 192 392 203
rect 384 180 385 182
rect 387 180 388 182
rect 384 174 388 180
rect 419 206 423 211
rect 475 211 476 213
rect 478 211 479 213
rect 475 209 479 211
rect 508 211 510 213
rect 512 211 514 213
rect 508 210 514 211
rect 539 211 540 213
rect 542 211 543 213
rect 539 209 543 211
rect 572 211 574 213
rect 576 211 578 213
rect 572 210 578 211
rect 603 211 604 213
rect 606 211 607 213
rect 603 209 607 211
rect 636 211 638 213
rect 640 211 642 213
rect 636 210 642 211
rect 419 204 420 206
rect 422 204 423 206
rect 419 202 423 204
rect 427 207 460 208
rect 427 205 456 207
rect 458 205 460 207
rect 427 204 460 205
rect 427 193 431 204
rect 408 192 431 193
rect 408 190 410 192
rect 412 190 431 192
rect 408 189 431 190
rect 408 183 412 189
rect 370 173 388 174
rect 370 171 372 173
rect 374 171 388 173
rect 370 170 388 171
rect 401 179 412 183
rect 401 173 405 179
rect 427 183 431 189
rect 435 199 439 201
rect 491 203 504 204
rect 491 201 493 203
rect 495 201 504 203
rect 491 200 504 201
rect 435 197 436 199
rect 438 197 439 199
rect 435 192 439 197
rect 500 196 516 200
rect 435 190 436 192
rect 438 191 439 192
rect 438 190 451 191
rect 435 187 451 190
rect 447 185 451 187
rect 447 183 452 185
rect 427 182 443 183
rect 427 180 439 182
rect 441 180 443 182
rect 427 179 443 180
rect 447 181 449 183
rect 451 181 452 183
rect 447 179 452 181
rect 401 171 402 173
rect 404 171 405 173
rect 401 169 405 171
rect 447 175 451 179
rect 427 171 451 175
rect 488 192 492 194
rect 320 166 340 167
rect 285 164 289 166
rect 296 165 302 166
rect 296 163 298 165
rect 300 163 302 165
rect 320 164 322 166
rect 324 164 340 166
rect 320 163 340 164
rect 427 168 431 171
rect 427 166 428 168
rect 430 166 431 168
rect 205 157 211 163
rect 296 157 302 163
rect 414 165 420 166
rect 414 163 416 165
rect 418 163 420 165
rect 427 164 431 166
rect 464 191 489 192
rect 464 189 466 191
rect 468 190 489 191
rect 491 190 492 192
rect 468 189 492 190
rect 464 188 492 189
rect 464 168 468 188
rect 488 178 492 188
rect 508 183 509 189
rect 512 179 516 196
rect 488 176 499 178
rect 488 174 496 176
rect 498 174 499 176
rect 512 177 517 179
rect 512 175 514 177
rect 516 175 517 177
rect 488 172 499 174
rect 502 173 517 175
rect 502 171 516 173
rect 464 167 470 168
rect 464 165 466 167
rect 468 165 470 167
rect 464 164 470 165
rect 474 167 480 168
rect 474 165 476 167
rect 478 165 480 167
rect 502 166 506 171
rect 555 203 568 204
rect 555 201 557 203
rect 559 201 568 203
rect 555 200 568 201
rect 564 196 580 200
rect 552 192 556 194
rect 360 160 366 161
rect 360 158 362 160
rect 364 158 366 160
rect 360 157 366 158
rect 379 160 385 161
rect 379 158 381 160
rect 383 158 385 160
rect 379 157 385 158
rect 414 157 420 163
rect 474 157 480 165
rect 491 165 506 166
rect 491 163 493 165
rect 495 163 506 165
rect 491 162 506 163
rect 509 165 513 167
rect 509 163 510 165
rect 512 163 513 165
rect 528 191 553 192
rect 528 189 530 191
rect 532 190 553 191
rect 555 190 556 192
rect 532 189 556 190
rect 528 188 556 189
rect 528 168 532 188
rect 552 178 556 188
rect 572 183 573 189
rect 576 179 580 196
rect 552 176 563 178
rect 552 174 560 176
rect 562 174 563 176
rect 576 177 581 179
rect 576 175 578 177
rect 580 175 581 177
rect 552 172 563 174
rect 566 173 581 175
rect 619 203 632 204
rect 619 201 621 203
rect 623 201 632 203
rect 619 200 632 201
rect 628 196 644 200
rect 616 192 620 194
rect 566 171 580 173
rect 528 167 534 168
rect 528 165 530 167
rect 532 165 534 167
rect 528 164 534 165
rect 538 167 544 168
rect 538 165 540 167
rect 542 165 544 167
rect 566 166 570 171
rect 509 157 513 163
rect 538 157 544 165
rect 555 165 570 166
rect 555 163 557 165
rect 559 163 570 165
rect 555 162 570 163
rect 573 165 577 167
rect 573 163 574 165
rect 576 163 577 165
rect 592 191 617 192
rect 592 189 594 191
rect 596 190 617 191
rect 619 190 620 192
rect 596 189 620 190
rect 592 188 620 189
rect 592 168 596 188
rect 616 178 620 188
rect 636 183 637 189
rect 640 179 644 196
rect 616 176 627 178
rect 616 174 624 176
rect 626 174 627 176
rect 640 177 645 179
rect 640 175 642 177
rect 644 175 645 177
rect 616 172 627 174
rect 630 173 645 175
rect 630 171 644 173
rect 592 167 598 168
rect 592 165 594 167
rect 596 165 598 167
rect 592 164 598 165
rect 602 167 608 168
rect 602 165 604 167
rect 606 165 608 167
rect 630 166 634 171
rect 573 157 577 163
rect 602 157 608 165
rect 619 165 634 166
rect 619 163 621 165
rect 623 163 634 165
rect 619 162 634 163
rect 637 165 641 167
rect 637 163 638 165
rect 640 163 641 165
rect 637 157 641 163
rect 47 135 53 141
rect 36 132 40 134
rect 47 133 49 135
rect 51 133 53 135
rect 47 132 53 133
rect 71 134 91 135
rect 71 132 73 134
rect 75 132 91 134
rect 36 130 37 132
rect 39 130 40 132
rect 71 131 91 132
rect 36 127 40 130
rect 16 123 40 127
rect 16 119 20 123
rect 62 127 66 129
rect 62 125 63 127
rect 65 125 66 127
rect 15 117 20 119
rect 15 115 16 117
rect 18 115 20 117
rect 24 118 40 119
rect 24 116 26 118
rect 28 116 40 118
rect 24 115 40 116
rect 15 113 20 115
rect 16 111 20 113
rect 16 108 32 111
rect 16 107 29 108
rect 28 106 29 107
rect 31 106 32 108
rect 28 101 32 106
rect 28 99 29 101
rect 31 99 32 101
rect 28 97 32 99
rect 36 109 40 115
rect 62 119 66 125
rect 55 115 66 119
rect 87 127 91 131
rect 151 135 157 141
rect 215 140 221 141
rect 215 138 217 140
rect 219 138 221 140
rect 215 137 221 138
rect 234 140 240 141
rect 234 138 236 140
rect 238 138 240 140
rect 234 137 240 138
rect 102 128 103 130
rect 87 123 99 127
rect 95 118 99 123
rect 95 116 96 118
rect 98 116 99 118
rect 55 109 59 115
rect 36 108 59 109
rect 36 106 55 108
rect 57 106 59 108
rect 36 105 59 106
rect 36 94 40 105
rect 95 104 99 116
rect 82 101 99 104
rect 82 99 83 101
rect 85 100 99 101
rect 85 99 86 100
rect 7 93 40 94
rect 7 91 9 93
rect 11 91 40 93
rect 7 90 40 91
rect 44 94 48 96
rect 44 92 45 94
rect 47 92 48 94
rect 44 87 48 92
rect 71 94 77 95
rect 71 92 73 94
rect 75 92 77 94
rect 44 85 45 87
rect 47 85 48 87
rect 71 85 77 92
rect 82 94 86 99
rect 140 132 144 134
rect 151 133 153 135
rect 155 133 157 135
rect 151 132 157 133
rect 175 134 195 135
rect 175 132 177 134
rect 179 132 195 134
rect 140 130 141 132
rect 143 130 144 132
rect 175 131 195 132
rect 140 127 144 130
rect 120 123 144 127
rect 120 119 124 123
rect 166 127 170 129
rect 166 125 167 127
rect 169 125 170 127
rect 119 117 124 119
rect 119 115 120 117
rect 122 115 124 117
rect 128 118 144 119
rect 128 116 130 118
rect 132 116 144 118
rect 128 115 144 116
rect 119 113 124 115
rect 120 111 124 113
rect 120 108 136 111
rect 120 107 133 108
rect 132 106 133 107
rect 135 106 136 108
rect 132 101 136 106
rect 132 99 133 101
rect 135 99 136 101
rect 132 97 136 99
rect 140 109 144 115
rect 166 119 170 125
rect 159 115 170 119
rect 191 127 195 131
rect 296 135 302 141
rect 360 140 366 141
rect 360 138 362 140
rect 364 138 366 140
rect 360 137 366 138
rect 379 140 385 141
rect 379 138 381 140
rect 383 138 385 140
rect 379 137 385 138
rect 206 128 207 130
rect 191 123 203 127
rect 199 118 203 123
rect 199 116 200 118
rect 202 116 203 118
rect 159 109 163 115
rect 140 108 163 109
rect 140 106 159 108
rect 161 106 163 108
rect 140 105 163 106
rect 82 92 83 94
rect 85 92 86 94
rect 82 90 86 92
rect 91 96 97 97
rect 91 94 93 96
rect 95 94 97 96
rect 140 94 144 105
rect 199 104 203 116
rect 285 132 289 134
rect 296 133 298 135
rect 300 133 302 135
rect 296 132 302 133
rect 320 134 340 135
rect 320 132 322 134
rect 324 132 340 134
rect 225 127 243 128
rect 225 125 227 127
rect 229 125 243 127
rect 225 124 243 125
rect 239 118 243 124
rect 239 116 240 118
rect 242 116 243 118
rect 218 111 224 112
rect 186 101 203 104
rect 186 99 187 101
rect 189 100 203 101
rect 189 99 190 100
rect 91 85 97 94
rect 111 93 144 94
rect 111 91 113 93
rect 115 91 144 93
rect 111 90 144 91
rect 148 94 152 96
rect 148 92 149 94
rect 151 92 152 94
rect 148 87 152 92
rect 175 94 181 95
rect 175 92 177 94
rect 179 92 181 94
rect 148 85 149 87
rect 151 85 152 87
rect 175 85 181 92
rect 186 94 190 99
rect 239 103 243 116
rect 228 99 243 103
rect 186 92 187 94
rect 189 92 190 94
rect 186 90 190 92
rect 195 96 201 97
rect 195 94 197 96
rect 199 94 201 96
rect 228 95 232 99
rect 246 95 247 106
rect 285 130 286 132
rect 288 130 289 132
rect 320 131 340 132
rect 285 127 289 130
rect 265 123 289 127
rect 265 119 269 123
rect 311 127 315 129
rect 311 125 312 127
rect 314 125 315 127
rect 264 117 269 119
rect 264 115 265 117
rect 267 115 269 117
rect 273 118 289 119
rect 273 116 275 118
rect 277 116 289 118
rect 273 115 289 116
rect 264 113 269 115
rect 265 111 269 113
rect 265 108 281 111
rect 265 107 278 108
rect 277 106 278 107
rect 280 106 281 108
rect 277 101 281 106
rect 277 99 278 101
rect 280 99 281 101
rect 277 97 281 99
rect 285 109 289 115
rect 311 119 315 125
rect 304 115 315 119
rect 336 127 340 131
rect 414 135 420 141
rect 414 133 416 135
rect 418 133 420 135
rect 414 132 420 133
rect 427 132 431 134
rect 351 128 352 130
rect 336 123 348 127
rect 344 118 348 123
rect 344 116 345 118
rect 347 116 348 118
rect 304 109 308 115
rect 285 108 308 109
rect 285 106 304 108
rect 306 106 308 108
rect 285 105 308 106
rect 195 85 201 94
rect 215 94 232 95
rect 215 92 217 94
rect 219 92 232 94
rect 215 91 232 92
rect 285 94 289 105
rect 344 104 348 116
rect 427 130 428 132
rect 430 130 431 132
rect 370 127 388 128
rect 370 125 372 127
rect 374 125 388 127
rect 370 124 388 125
rect 384 118 388 124
rect 384 116 385 118
rect 387 116 388 118
rect 363 111 369 112
rect 331 101 348 104
rect 331 99 332 101
rect 334 100 348 101
rect 334 99 335 100
rect 256 93 289 94
rect 256 91 258 93
rect 260 91 289 93
rect 256 90 289 91
rect 293 94 297 96
rect 293 92 294 94
rect 296 92 297 94
rect 234 87 240 88
rect 234 85 236 87
rect 238 85 240 87
rect 293 87 297 92
rect 320 94 326 95
rect 320 92 322 94
rect 324 92 326 94
rect 293 85 294 87
rect 296 85 297 87
rect 320 85 326 92
rect 331 94 335 99
rect 384 103 388 116
rect 401 127 405 129
rect 401 125 402 127
rect 404 125 405 127
rect 401 119 405 125
rect 427 127 431 130
rect 427 123 451 127
rect 401 115 412 119
rect 373 99 388 103
rect 331 92 332 94
rect 334 92 335 94
rect 331 90 335 92
rect 340 96 346 97
rect 340 94 342 96
rect 344 94 346 96
rect 373 95 377 99
rect 391 95 392 106
rect 340 85 346 94
rect 360 94 377 95
rect 360 92 362 94
rect 364 92 377 94
rect 360 91 377 92
rect 408 109 412 115
rect 447 119 451 123
rect 427 118 443 119
rect 427 116 439 118
rect 441 116 443 118
rect 427 115 443 116
rect 447 117 452 119
rect 447 115 449 117
rect 451 115 452 117
rect 427 109 431 115
rect 447 113 452 115
rect 447 111 451 113
rect 408 108 431 109
rect 408 106 410 108
rect 412 106 431 108
rect 408 105 431 106
rect 419 94 423 96
rect 419 92 420 94
rect 422 92 423 94
rect 379 87 385 88
rect 379 85 381 87
rect 383 85 385 87
rect 419 87 423 92
rect 427 94 431 105
rect 435 108 451 111
rect 435 106 436 108
rect 438 107 451 108
rect 438 106 439 107
rect 435 101 439 106
rect 464 133 470 134
rect 464 131 466 133
rect 468 131 470 133
rect 464 130 470 131
rect 474 133 480 141
rect 474 131 476 133
rect 478 131 480 133
rect 491 135 506 136
rect 491 133 493 135
rect 495 133 506 135
rect 491 132 506 133
rect 474 130 480 131
rect 464 110 468 130
rect 502 127 506 132
rect 509 135 513 141
rect 509 133 510 135
rect 512 133 513 135
rect 509 131 513 133
rect 488 124 499 126
rect 488 122 496 124
rect 498 122 499 124
rect 502 125 516 127
rect 502 123 517 125
rect 488 120 499 122
rect 512 121 514 123
rect 516 121 517 123
rect 488 110 492 120
rect 512 119 517 121
rect 464 109 492 110
rect 464 107 466 109
rect 468 108 492 109
rect 468 107 489 108
rect 464 106 489 107
rect 491 106 492 108
rect 508 109 509 115
rect 488 104 492 106
rect 435 99 436 101
rect 438 99 439 101
rect 435 97 439 99
rect 512 102 516 119
rect 500 98 516 102
rect 528 133 534 134
rect 528 131 530 133
rect 532 131 534 133
rect 528 130 534 131
rect 538 133 544 141
rect 538 131 540 133
rect 542 131 544 133
rect 555 135 570 136
rect 555 133 557 135
rect 559 133 570 135
rect 555 132 570 133
rect 538 130 544 131
rect 528 110 532 130
rect 566 127 570 132
rect 573 135 577 141
rect 573 133 574 135
rect 576 133 577 135
rect 573 131 577 133
rect 552 124 563 126
rect 552 122 560 124
rect 562 122 563 124
rect 566 125 580 127
rect 566 123 581 125
rect 552 120 563 122
rect 576 121 578 123
rect 580 121 581 123
rect 552 110 556 120
rect 576 119 581 121
rect 528 109 556 110
rect 528 107 530 109
rect 532 108 556 109
rect 532 107 553 108
rect 528 106 553 107
rect 555 106 556 108
rect 572 109 573 115
rect 552 104 556 106
rect 427 93 460 94
rect 427 91 456 93
rect 458 91 460 93
rect 427 90 460 91
rect 491 97 504 98
rect 491 95 493 97
rect 495 95 504 97
rect 491 94 504 95
rect 576 102 580 119
rect 564 98 580 102
rect 555 97 568 98
rect 555 95 557 97
rect 559 95 568 97
rect 592 133 598 134
rect 592 131 594 133
rect 596 131 598 133
rect 592 130 598 131
rect 602 133 608 141
rect 602 131 604 133
rect 606 131 608 133
rect 619 135 634 136
rect 619 133 621 135
rect 623 133 634 135
rect 619 132 634 133
rect 602 130 608 131
rect 592 110 596 130
rect 630 127 634 132
rect 637 135 641 141
rect 637 133 638 135
rect 640 133 641 135
rect 637 131 641 133
rect 616 124 627 126
rect 616 122 624 124
rect 626 122 627 124
rect 630 125 644 127
rect 630 123 645 125
rect 616 120 627 122
rect 640 121 642 123
rect 644 121 645 123
rect 616 110 620 120
rect 640 119 645 121
rect 592 109 620 110
rect 592 107 594 109
rect 596 108 620 109
rect 596 107 617 108
rect 592 106 617 107
rect 619 106 620 108
rect 636 109 637 115
rect 616 104 620 106
rect 555 94 568 95
rect 640 102 644 119
rect 628 98 644 102
rect 619 97 632 98
rect 619 95 621 97
rect 623 95 632 97
rect 619 94 632 95
rect 419 85 420 87
rect 422 85 423 87
rect 475 87 479 89
rect 475 85 476 87
rect 478 85 479 87
rect 508 87 514 88
rect 508 85 510 87
rect 512 85 514 87
rect 539 87 543 89
rect 539 85 540 87
rect 542 85 543 87
rect 572 87 578 88
rect 572 85 574 87
rect 576 85 578 87
rect 603 87 607 89
rect 603 85 604 87
rect 606 85 607 87
rect 636 87 642 88
rect 636 85 638 87
rect 640 85 642 87
rect 18 67 20 69
rect 22 67 24 69
rect 18 66 24 67
rect 26 62 43 63
rect 26 60 39 62
rect 41 60 43 62
rect 26 59 43 60
rect 57 60 63 69
rect 11 48 12 59
rect 26 55 30 59
rect 57 58 59 60
rect 61 58 63 60
rect 57 57 63 58
rect 68 62 72 64
rect 68 60 69 62
rect 71 60 72 62
rect 15 51 30 55
rect 15 38 19 51
rect 68 55 72 60
rect 77 62 83 69
rect 106 67 107 69
rect 109 67 110 69
rect 77 60 79 62
rect 81 60 83 62
rect 77 59 83 60
rect 106 62 110 67
rect 106 60 107 62
rect 109 60 110 62
rect 106 58 110 60
rect 114 63 147 64
rect 114 61 143 63
rect 145 61 147 63
rect 114 60 147 61
rect 161 60 167 69
rect 68 54 69 55
rect 55 53 69 54
rect 71 53 72 55
rect 55 50 72 53
rect 34 42 40 43
rect 15 36 16 38
rect 18 36 19 38
rect 15 30 19 36
rect 15 29 33 30
rect 15 27 29 29
rect 31 27 33 29
rect 15 26 33 27
rect 55 38 59 50
rect 114 49 118 60
rect 161 58 163 60
rect 165 58 167 60
rect 161 57 167 58
rect 172 62 176 64
rect 172 60 173 62
rect 175 60 176 62
rect 95 48 118 49
rect 95 46 97 48
rect 99 46 118 48
rect 95 45 118 46
rect 95 39 99 45
rect 55 36 56 38
rect 58 36 59 38
rect 55 31 59 36
rect 55 27 67 31
rect 51 24 52 26
rect 63 23 67 27
rect 88 35 99 39
rect 88 29 92 35
rect 114 39 118 45
rect 122 55 126 57
rect 122 53 123 55
rect 125 53 126 55
rect 122 48 126 53
rect 122 46 123 48
rect 125 47 126 48
rect 125 46 138 47
rect 122 43 138 46
rect 134 41 138 43
rect 134 39 139 41
rect 114 38 130 39
rect 114 36 126 38
rect 128 36 130 38
rect 114 35 130 36
rect 134 37 136 39
rect 138 37 139 39
rect 134 35 139 37
rect 88 27 89 29
rect 91 27 92 29
rect 88 25 92 27
rect 134 31 138 35
rect 114 27 138 31
rect 114 24 118 27
rect 63 22 83 23
rect 114 22 115 24
rect 117 22 118 24
rect 63 20 79 22
rect 81 20 83 22
rect 63 19 83 20
rect 101 21 107 22
rect 101 19 103 21
rect 105 19 107 21
rect 114 20 118 22
rect 172 55 176 60
rect 181 62 187 69
rect 210 67 211 69
rect 213 67 214 69
rect 181 60 183 62
rect 185 60 187 62
rect 181 59 187 60
rect 210 62 214 67
rect 293 67 294 69
rect 296 67 297 69
rect 210 60 211 62
rect 213 60 214 62
rect 210 58 214 60
rect 218 63 251 64
rect 218 61 247 63
rect 249 61 251 63
rect 218 60 251 61
rect 256 63 289 64
rect 256 61 258 63
rect 260 61 289 63
rect 256 60 289 61
rect 172 54 173 55
rect 159 53 173 54
rect 175 53 176 55
rect 159 50 176 53
rect 159 38 163 50
rect 218 49 222 60
rect 199 48 222 49
rect 199 46 201 48
rect 203 46 222 48
rect 199 45 222 46
rect 199 39 203 45
rect 159 36 160 38
rect 162 36 163 38
rect 159 31 163 36
rect 159 27 171 31
rect 155 24 156 26
rect 18 16 24 17
rect 18 14 20 16
rect 22 14 24 16
rect 18 13 24 14
rect 37 16 43 17
rect 37 14 39 16
rect 41 14 43 16
rect 37 13 43 14
rect 101 13 107 19
rect 167 23 171 27
rect 192 35 203 39
rect 192 29 196 35
rect 218 39 222 45
rect 226 55 230 57
rect 226 53 227 55
rect 229 53 230 55
rect 226 48 230 53
rect 226 46 227 48
rect 229 47 230 48
rect 229 46 242 47
rect 226 43 242 46
rect 238 41 242 43
rect 238 39 243 41
rect 218 38 234 39
rect 218 36 230 38
rect 232 36 234 38
rect 218 35 234 36
rect 238 37 240 39
rect 242 37 243 39
rect 238 35 243 37
rect 192 27 193 29
rect 195 27 196 29
rect 192 25 196 27
rect 238 31 242 35
rect 218 27 242 31
rect 218 24 222 27
rect 167 22 187 23
rect 218 22 219 24
rect 221 22 222 24
rect 167 20 183 22
rect 185 20 187 22
rect 167 19 187 20
rect 205 21 211 22
rect 205 19 207 21
rect 209 19 211 21
rect 218 20 222 22
rect 277 55 281 57
rect 277 53 278 55
rect 280 53 281 55
rect 277 48 281 53
rect 277 47 278 48
rect 265 46 278 47
rect 280 46 281 48
rect 265 43 281 46
rect 285 49 289 60
rect 293 62 297 67
rect 293 60 294 62
rect 296 60 297 62
rect 293 58 297 60
rect 320 62 326 69
rect 320 60 322 62
rect 324 60 326 62
rect 320 59 326 60
rect 331 62 335 64
rect 331 60 332 62
rect 334 60 335 62
rect 285 48 308 49
rect 285 46 304 48
rect 306 46 308 48
rect 285 45 308 46
rect 265 41 269 43
rect 264 39 269 41
rect 285 39 289 45
rect 264 37 265 39
rect 267 37 269 39
rect 264 35 269 37
rect 273 38 289 39
rect 273 36 275 38
rect 277 36 289 38
rect 273 35 289 36
rect 265 31 269 35
rect 304 39 308 45
rect 331 55 335 60
rect 340 60 346 69
rect 379 67 381 69
rect 383 67 385 69
rect 379 66 385 67
rect 419 67 420 69
rect 422 67 423 69
rect 340 58 342 60
rect 344 58 346 60
rect 360 62 377 63
rect 360 60 362 62
rect 364 60 377 62
rect 360 59 377 60
rect 340 57 346 58
rect 331 53 332 55
rect 334 54 335 55
rect 334 53 348 54
rect 331 50 348 53
rect 304 35 315 39
rect 265 27 289 31
rect 285 24 289 27
rect 311 29 315 35
rect 311 27 312 29
rect 314 27 315 29
rect 311 25 315 27
rect 344 38 348 50
rect 344 36 345 38
rect 347 36 348 38
rect 344 31 348 36
rect 336 27 348 31
rect 285 22 286 24
rect 288 22 289 24
rect 336 23 340 27
rect 351 24 352 26
rect 373 55 377 59
rect 373 51 388 55
rect 363 42 369 43
rect 384 38 388 51
rect 391 48 392 59
rect 384 36 385 38
rect 387 36 388 38
rect 384 30 388 36
rect 419 62 423 67
rect 475 67 476 69
rect 478 67 479 69
rect 475 65 479 67
rect 508 67 510 69
rect 512 67 514 69
rect 508 66 514 67
rect 539 67 540 69
rect 542 67 543 69
rect 539 65 543 67
rect 572 67 574 69
rect 576 67 578 69
rect 572 66 578 67
rect 603 67 604 69
rect 606 67 607 69
rect 603 65 607 67
rect 636 67 638 69
rect 640 67 642 69
rect 636 66 642 67
rect 419 60 420 62
rect 422 60 423 62
rect 419 58 423 60
rect 427 63 460 64
rect 427 61 456 63
rect 458 61 460 63
rect 427 60 460 61
rect 427 49 431 60
rect 408 48 431 49
rect 408 46 410 48
rect 412 46 431 48
rect 408 45 431 46
rect 408 39 412 45
rect 370 29 388 30
rect 370 27 372 29
rect 374 27 388 29
rect 370 26 388 27
rect 401 35 412 39
rect 401 29 405 35
rect 427 39 431 45
rect 435 55 439 57
rect 491 59 504 60
rect 491 57 493 59
rect 495 57 504 59
rect 491 56 504 57
rect 435 53 436 55
rect 438 53 439 55
rect 435 48 439 53
rect 500 52 516 56
rect 435 46 436 48
rect 438 47 439 48
rect 438 46 451 47
rect 435 43 451 46
rect 447 41 451 43
rect 447 39 452 41
rect 427 38 443 39
rect 427 36 439 38
rect 441 36 443 38
rect 427 35 443 36
rect 447 37 449 39
rect 451 37 452 39
rect 447 35 452 37
rect 401 27 402 29
rect 404 27 405 29
rect 401 25 405 27
rect 447 31 451 35
rect 427 27 451 31
rect 488 48 492 50
rect 320 22 340 23
rect 285 20 289 22
rect 296 21 302 22
rect 296 19 298 21
rect 300 19 302 21
rect 320 20 322 22
rect 324 20 340 22
rect 320 19 340 20
rect 427 24 431 27
rect 427 22 428 24
rect 430 22 431 24
rect 205 13 211 19
rect 296 13 302 19
rect 414 21 420 22
rect 414 19 416 21
rect 418 19 420 21
rect 427 20 431 22
rect 464 47 489 48
rect 464 45 466 47
rect 468 46 489 47
rect 491 46 492 48
rect 468 45 492 46
rect 464 44 492 45
rect 464 24 468 44
rect 488 34 492 44
rect 508 39 509 45
rect 512 35 516 52
rect 488 32 499 34
rect 488 30 496 32
rect 498 30 499 32
rect 512 33 517 35
rect 512 31 514 33
rect 516 31 517 33
rect 488 28 499 30
rect 502 29 517 31
rect 502 27 516 29
rect 464 23 470 24
rect 464 21 466 23
rect 468 21 470 23
rect 464 20 470 21
rect 474 23 480 24
rect 474 21 476 23
rect 478 21 480 23
rect 502 22 506 27
rect 555 59 568 60
rect 555 57 557 59
rect 559 57 568 59
rect 555 56 568 57
rect 564 52 580 56
rect 552 48 556 50
rect 360 16 366 17
rect 360 14 362 16
rect 364 14 366 16
rect 360 13 366 14
rect 379 16 385 17
rect 379 14 381 16
rect 383 14 385 16
rect 379 13 385 14
rect 414 13 420 19
rect 474 13 480 21
rect 491 21 506 22
rect 491 19 493 21
rect 495 19 506 21
rect 491 18 506 19
rect 509 21 513 23
rect 509 19 510 21
rect 512 19 513 21
rect 528 47 553 48
rect 528 45 530 47
rect 532 46 553 47
rect 555 46 556 48
rect 532 45 556 46
rect 528 44 556 45
rect 528 24 532 44
rect 552 34 556 44
rect 572 39 573 45
rect 576 35 580 52
rect 552 32 563 34
rect 552 30 560 32
rect 562 30 563 32
rect 576 33 581 35
rect 576 31 578 33
rect 580 31 581 33
rect 552 28 563 30
rect 566 29 581 31
rect 619 59 632 60
rect 619 57 621 59
rect 623 57 632 59
rect 619 56 632 57
rect 628 52 644 56
rect 616 48 620 50
rect 566 27 580 29
rect 528 23 534 24
rect 528 21 530 23
rect 532 21 534 23
rect 528 20 534 21
rect 538 23 544 24
rect 538 21 540 23
rect 542 21 544 23
rect 566 22 570 27
rect 509 13 513 19
rect 538 13 544 21
rect 555 21 570 22
rect 555 19 557 21
rect 559 19 570 21
rect 555 18 570 19
rect 573 21 577 23
rect 573 19 574 21
rect 576 19 577 21
rect 592 47 617 48
rect 592 45 594 47
rect 596 46 617 47
rect 619 46 620 48
rect 596 45 620 46
rect 592 44 620 45
rect 592 24 596 44
rect 616 34 620 44
rect 636 39 637 45
rect 640 35 644 52
rect 616 32 627 34
rect 616 30 624 32
rect 626 30 627 32
rect 640 33 645 35
rect 640 31 642 33
rect 644 31 645 33
rect 616 28 627 30
rect 630 29 645 31
rect 630 27 644 29
rect 592 23 598 24
rect 592 21 594 23
rect 596 21 598 23
rect 592 20 598 21
rect 602 23 608 24
rect 602 21 604 23
rect 606 21 608 23
rect 630 22 634 27
rect 573 13 577 19
rect 602 13 608 21
rect 619 21 634 22
rect 619 19 621 21
rect 623 19 634 21
rect 619 18 634 19
rect 637 21 641 23
rect 637 19 638 21
rect 640 19 641 21
rect 637 13 641 19
<< via1 >>
rect 4 576 6 578
rect 55 557 57 559
rect 19 531 21 533
rect 80 557 82 559
rect 89 548 91 550
rect 63 533 65 535
rect 81 540 83 542
rect 104 548 106 550
rect 72 533 74 535
rect 159 557 161 559
rect 112 540 114 542
rect 184 557 186 559
rect 167 533 169 535
rect 216 548 218 550
rect 176 533 178 535
rect 208 535 210 537
rect 216 535 218 537
rect 303 556 305 558
rect 257 531 259 533
rect 329 556 331 558
rect 353 565 355 567
rect 313 532 315 534
rect 361 556 363 558
rect 321 532 323 534
rect 411 556 413 558
rect 393 541 395 543
rect 361 531 363 533
rect 457 556 459 558
rect 402 531 404 533
rect 472 556 474 558
rect 497 541 499 543
rect 536 556 538 558
rect 585 556 587 558
rect 561 541 563 543
rect 521 532 523 534
rect 466 523 468 525
rect 600 556 602 558
rect 625 539 627 541
rect 530 523 532 525
rect 594 523 596 525
rect 252 503 254 505
rect 8 470 10 472
rect 40 481 42 483
rect 48 481 50 483
rect 80 483 82 485
rect 40 468 42 470
rect 89 483 91 485
rect 72 459 74 461
rect 144 476 146 478
rect 97 459 99 461
rect 184 483 186 485
rect 152 468 154 470
rect 175 476 177 478
rect 193 483 195 485
rect 177 468 179 470
rect 176 459 178 461
rect 243 484 245 486
rect 201 459 203 461
rect 257 484 259 486
rect 313 485 315 487
rect 321 485 323 487
rect 303 460 305 462
rect 329 459 331 461
rect 361 485 363 487
rect 393 475 395 477
rect 465 493 467 495
rect 402 485 404 487
rect 361 459 363 461
rect 411 459 413 461
rect 457 460 459 462
rect 353 451 355 453
rect 472 460 474 462
rect 497 475 499 477
rect 521 484 523 486
rect 530 493 532 495
rect 536 460 538 462
rect 561 475 563 477
rect 594 493 596 495
rect 585 460 587 462
rect 600 460 602 462
rect 625 477 627 479
rect 4 442 6 444
rect 4 432 6 434
rect 55 413 57 415
rect 19 387 21 389
rect 80 413 82 415
rect 81 404 83 406
rect 63 389 65 391
rect 81 396 83 398
rect 104 404 106 406
rect 72 389 74 391
rect 159 413 161 415
rect 112 396 114 398
rect 184 413 186 415
rect 167 389 169 391
rect 216 404 218 406
rect 176 389 178 391
rect 208 391 210 393
rect 216 391 218 393
rect 248 407 250 409
rect 303 412 305 414
rect 257 387 259 389
rect 329 412 331 414
rect 353 421 355 423
rect 312 387 314 389
rect 361 412 363 414
rect 321 387 323 389
rect 412 412 414 414
rect 393 397 395 399
rect 361 387 363 389
rect 457 412 459 414
rect 401 387 403 389
rect 472 412 474 414
rect 497 397 499 399
rect 536 412 538 414
rect 585 412 587 414
rect 561 396 563 398
rect 521 388 523 390
rect 465 379 467 381
rect 600 412 602 414
rect 625 395 627 397
rect 530 379 532 381
rect 594 379 596 381
rect 252 368 254 370
rect 252 359 254 361
rect 8 324 10 326
rect 40 337 42 339
rect 48 337 50 339
rect 80 339 82 341
rect 40 324 42 326
rect 89 339 91 341
rect 72 315 74 317
rect 144 332 146 334
rect 97 315 99 317
rect 184 339 186 341
rect 152 324 154 326
rect 175 332 177 334
rect 193 339 195 341
rect 176 315 178 317
rect 237 341 239 343
rect 201 315 203 317
rect 257 340 259 342
rect 312 340 314 342
rect 321 340 323 342
rect 303 315 305 317
rect 329 316 331 318
rect 361 340 363 342
rect 393 331 395 333
rect 465 349 467 351
rect 401 340 403 342
rect 361 315 363 317
rect 413 316 415 318
rect 457 316 459 318
rect 353 307 355 309
rect 472 316 474 318
rect 497 331 499 333
rect 521 340 523 342
rect 530 349 532 351
rect 536 316 538 318
rect 561 331 563 333
rect 594 349 596 351
rect 585 316 587 318
rect 600 316 602 318
rect 625 333 627 335
rect 4 296 6 298
rect 4 288 6 290
rect 55 269 57 271
rect 19 243 21 245
rect 80 269 82 271
rect 89 260 91 262
rect 63 245 65 247
rect 81 252 83 254
rect 104 260 106 262
rect 72 245 74 247
rect 159 269 161 271
rect 112 252 114 254
rect 184 269 186 271
rect 167 245 169 247
rect 216 260 218 262
rect 176 245 178 247
rect 208 247 210 249
rect 216 247 218 249
rect 248 257 250 259
rect 303 268 305 270
rect 257 243 259 245
rect 329 269 331 271
rect 353 277 355 279
rect 312 243 314 245
rect 361 268 363 270
rect 321 243 323 245
rect 412 269 414 271
rect 393 253 395 255
rect 361 243 363 245
rect 457 268 459 270
rect 401 243 403 245
rect 472 268 474 270
rect 497 253 499 255
rect 536 268 538 270
rect 585 268 587 270
rect 561 253 563 255
rect 521 244 523 246
rect 465 235 467 237
rect 600 268 602 270
rect 625 251 627 253
rect 529 235 531 237
rect 594 235 596 237
rect 252 225 254 227
rect 252 215 254 217
rect 8 182 10 184
rect 40 193 42 195
rect 48 193 50 195
rect 80 195 82 197
rect 40 180 42 182
rect 89 195 91 197
rect 72 171 74 173
rect 144 188 146 190
rect 97 171 99 173
rect 184 195 186 197
rect 152 180 154 182
rect 175 188 177 190
rect 193 195 195 197
rect 177 180 179 182
rect 176 171 178 173
rect 243 196 245 198
rect 201 171 203 173
rect 257 196 259 198
rect 312 196 314 198
rect 321 196 323 198
rect 303 172 305 174
rect 329 171 331 173
rect 361 196 363 198
rect 393 187 395 189
rect 465 205 467 207
rect 401 196 403 198
rect 361 171 363 173
rect 412 172 414 174
rect 457 172 459 174
rect 353 163 355 165
rect 472 172 474 174
rect 497 187 499 189
rect 521 196 523 198
rect 529 205 531 207
rect 536 172 538 174
rect 561 187 563 189
rect 594 205 596 207
rect 585 172 587 174
rect 600 172 602 174
rect 625 189 627 191
rect 4 154 6 156
rect 4 144 6 146
rect 55 125 57 127
rect 19 99 21 101
rect 80 125 82 127
rect 81 116 83 118
rect 63 101 65 103
rect 81 108 83 110
rect 104 116 106 118
rect 72 101 74 103
rect 159 125 161 127
rect 112 108 114 110
rect 184 125 186 127
rect 167 101 169 103
rect 216 116 218 118
rect 176 101 178 103
rect 208 103 210 105
rect 216 103 218 105
rect 248 118 250 120
rect 303 124 305 126
rect 257 99 259 101
rect 329 124 331 126
rect 353 133 355 135
rect 312 99 314 101
rect 361 125 363 127
rect 321 99 323 101
rect 412 125 414 127
rect 393 108 395 110
rect 361 99 363 101
rect 457 124 459 126
rect 401 99 403 101
rect 472 124 474 126
rect 497 108 499 110
rect 536 124 538 126
rect 585 124 587 126
rect 561 108 563 110
rect 521 100 523 102
rect 465 91 467 93
rect 600 124 602 126
rect 625 107 627 109
rect 529 91 531 93
rect 594 91 596 93
rect 252 80 254 82
rect 8 36 10 38
rect 40 49 42 51
rect 48 49 50 51
rect 80 51 82 53
rect 40 36 42 38
rect 89 51 91 53
rect 72 27 74 29
rect 144 44 146 46
rect 97 27 99 29
rect 184 51 186 53
rect 152 36 154 38
rect 175 44 177 46
rect 193 51 195 53
rect 176 27 178 29
rect 248 43 250 45
rect 201 27 203 29
rect 257 52 259 54
rect 312 52 314 54
rect 321 52 323 54
rect 303 27 305 29
rect 329 27 331 29
rect 361 53 363 55
rect 393 43 395 45
rect 465 61 467 63
rect 401 52 403 54
rect 361 27 363 29
rect 412 28 414 30
rect 457 28 459 30
rect 353 19 355 21
rect 478 28 480 30
rect 497 43 499 45
rect 521 52 523 54
rect 530 61 532 63
rect 536 28 538 30
rect 561 43 563 45
rect 594 61 596 63
rect 585 28 587 30
rect 600 28 602 30
rect 625 45 627 47
rect 4 8 6 10
<< via2 >>
rect 4 576 6 578
rect 184 557 186 559
rect 19 531 21 533
rect 252 503 254 505
rect 243 484 245 486
rect 97 459 99 461
rect 4 442 6 444
rect 4 432 6 434
rect 184 413 186 415
rect 329 556 331 558
rect 561 541 563 543
rect 466 523 468 525
rect 594 523 596 525
rect 465 493 467 495
rect 594 493 596 495
rect 561 475 563 477
rect 329 459 331 461
rect 19 387 21 389
rect 252 368 254 370
rect 252 359 254 361
rect 237 341 239 343
rect 329 412 331 414
rect 561 396 563 398
rect 465 379 467 381
rect 594 379 596 381
rect 465 349 467 351
rect 594 349 596 351
rect 561 331 563 333
rect 97 315 99 317
rect 329 316 331 318
rect 4 296 6 298
rect 4 288 6 290
rect 159 269 161 271
rect 19 243 21 245
rect 252 225 254 227
rect 252 215 254 217
rect 243 196 245 198
rect 97 171 99 173
rect 4 154 6 156
rect 4 144 6 146
rect 159 125 161 127
rect 329 269 331 271
rect 561 253 563 255
rect 465 235 467 237
rect 594 235 596 237
rect 465 205 467 207
rect 594 205 596 207
rect 561 187 563 189
rect 329 171 331 173
rect 19 99 21 101
rect 252 80 254 82
rect 248 43 250 45
rect 329 124 331 126
rect 561 108 563 110
rect 465 91 467 93
rect 594 91 596 93
rect 465 61 467 63
rect 594 61 596 63
rect 561 43 563 45
rect 4 8 6 10
<< via3 >>
rect 184 557 186 559
rect 329 556 331 558
rect 561 541 563 543
rect 19 531 21 533
rect 243 484 245 486
rect 97 459 99 461
rect 184 413 186 415
rect 19 387 21 389
rect 329 459 331 461
rect 329 412 331 414
rect 561 475 563 477
rect 561 396 563 398
rect 237 341 239 343
rect 97 315 99 317
rect 159 269 161 271
rect 19 243 21 245
rect 329 316 331 318
rect 329 269 331 271
rect 561 331 563 333
rect 561 253 563 255
rect 243 196 245 198
rect 97 171 99 173
rect 159 125 161 127
rect 19 99 21 101
rect 329 171 331 173
rect 329 124 331 126
rect 561 187 563 189
rect 561 108 563 110
<< labels >>
rlabel alu0 90 32 90 32 6 bn
rlabel alu0 136 37 136 37 6 an
rlabel alu0 57 40 57 40 6 zn
rlabel alu1 145 33 145 33 1 s
rlabel alu1 57 21 57 21 1 co
rlabel alu0 161 39 161 39 1 zn_1
rlabel alu0 194 32 194 32 1 bn_1
rlabel alu0 220 24 220 24 1 an_1
rlabel alu1 25 9 25 9 6 vss
rlabel alu1 161 21 161 21 1 c1
rlabel alu0 34 61 34 61 1 zn_2
rlabel alu1 9 41 9 41 1 cout0
rlabel alu1 249 32 249 32 1 sum0
rlabel alu1 37 81 37 81 2 vdd
rlabel alu1 9 121 9 121 1 sum1
rlabel alu0 38 130 38 130 1 1_an_1
rlabel alu0 64 122 64 122 1 1_bn_1
rlabel alu0 97 115 97 115 1 1_zn_1
rlabel alu1 97 132 97 132 1 1_c1
rlabel alu0 122 117 122 117 1 1_an
rlabel alu1 113 120 113 120 1 1_s
rlabel alu0 168 122 168 122 1 1_bn
rlabel alu0 201 114 201 114 1 1_zn
rlabel alu1 201 133 201 133 1 1_co
rlabel alu0 224 93 224 93 1 1_zn_2
rlabel alu1 249 113 249 113 1 cout1
rlabel alu1 9 184 9 184 1 cout2
rlabel alu0 34 205 34 205 1 2_zn_2
rlabel alu1 57 165 57 165 1 2_co
rlabel alu0 57 184 57 184 1 2_zn
rlabel alu0 90 176 90 176 1 2_bn
rlabel alu0 136 181 136 181 1 2_an
rlabel alu1 145 177 145 177 1 2_s
rlabel alu1 161 165 161 165 1 2_c1
rlabel alu0 161 183 161 183 1 2_zn_1
rlabel alu0 194 176 194 176 1 2_bn_1
rlabel alu0 220 168 220 168 1 2_an_1
rlabel alu1 249 177 249 177 1 sum2
rlabel alu1 37 289 37 289 2 vss
rlabel alu1 9 264 9 264 1 sum3
rlabel alu1 249 257 249 257 1 cout3
rlabel alu0 38 274 38 274 1 3_an_1
rlabel alu0 64 266 64 266 1 3_bn_1
rlabel alu0 97 259 97 259 1 3_zn_1
rlabel alu1 113 264 113 264 1 3_s
rlabel alu0 122 261 122 261 1 3_an
rlabel alu1 97 277 97 277 1 3_c1
rlabel alu0 168 266 168 266 1 3_bn
rlabel alu0 201 258 201 258 1 3_zn
rlabel alu1 201 277 201 277 1 3_co
rlabel alu0 224 237 224 237 1 3_zn_2
rlabel polyct1 105 33 105 33 1 A0
rlabel polyct1 153 121 153 121 1 A1
rlabel polyct1 105 177 105 177 1 A2
rlabel polyct1 153 265 153 265 1 A3
rlabel via1 81 53 81 53 1 tb0
rlabel via1 177 101 177 101 1 tb1
rlabel via1 81 197 81 197 1 tb2
rlabel alu2 177 244 177 244 1 tb3
rlabel alu1 286 9 286 9 4 vss
rlabel alu1 313 61 313 61 1 B0
rlabel polyct1 298 31 298 31 1 MODE
rlabel alu0 267 38 267 38 1 an_2
rlabel alu0 313 32 313 32 1 bn_2
rlabel alu1 313 94 313 94 1 B1
rlabel polyct1 298 121 298 121 1 MODE
rlabel alu0 267 116 267 116 1 1_an_2
rlabel alu0 273 92 273 92 1 1_bn_2
rlabel polyct1 298 177 298 177 1 MODE
rlabel alu1 313 205 313 205 1 B2
rlabel alu0 267 182 267 182 1 2_an_2
rlabel alu0 273 206 273 206 1 2_bn_2
rlabel alu1 286 289 286 289 2 vss
rlabel alu1 313 238 313 238 1 B3
rlabel polyct1 298 265 298 265 1 MODE
rlabel alu0 267 261 267 261 1 3_an_2
rlabel alu0 277 262 277 262 1 3_bn_2
rlabel alu1 25 297 25 297 6 vss
rlabel alu1 37 369 37 369 2 vdd
rlabel alu1 37 577 37 577 2 vss
rlabel alu1 37 513 37 513 2 vdd
rlabel alu1 286 297 286 297 4 vss
rlabel polyct1 298 319 298 319 1 MODE
rlabel polyct1 298 409 298 409 1 MODE
rlabel polyct1 298 465 298 465 1 MODE
rlabel alu1 286 577 286 577 2 vss
rlabel polyct1 298 553 298 553 1 MODE
rlabel alu1 9 329 9 329 1 cout4
rlabel alu0 34 349 34 349 1 4_zn_2
rlabel alu0 57 328 57 328 1 4_zn
rlabel alu1 57 309 57 309 1 4_co
rlabel via1 81 341 81 341 1 tb4
rlabel alu0 90 320 90 320 1 4_bn
rlabel polyct1 105 321 105 321 1 A4
rlabel alu0 136 325 136 325 1 4_an
rlabel alu1 145 321 145 321 1 4_s
rlabel alu1 161 309 161 309 1 4_c1
rlabel alu0 161 327 161 327 1 4_zn_1
rlabel alu0 194 320 194 320 1 4_bn_1
rlabel alu0 220 312 220 312 1 4_an_1
rlabel alu1 249 320 249 320 1 sum4
rlabel alu0 267 326 267 326 1 4_an_2
rlabel alu0 313 320 313 320 1 4_bn_2
rlabel alu1 313 349 313 349 1 B4
rlabel alu1 313 383 313 383 1 B5
rlabel alu0 273 380 273 380 1 5_bn_2
rlabel alu0 267 404 267 404 1 5_an_2
rlabel alu0 224 381 224 381 1 5_zn_2
rlabel alu1 201 421 201 421 1 5_co
rlabel alu0 201 402 201 402 1 5_zn
rlabel via1 177 389 177 389 1 tb5
rlabel alu0 168 410 168 410 1 5_bn
rlabel polyct1 153 409 153 409 1 A5
rlabel alu0 122 405 122 405 1 5_an
rlabel alu1 113 408 113 408 1 5_s
rlabel alu0 97 404 97 404 1 5_zn_1
rlabel alu1 97 420 97 420 1 5_c1
rlabel alu0 64 410 64 410 1 5_bn_1
rlabel alu0 38 418 38 418 1 5_an_1
rlabel alu1 9 410 9 410 1 sum5
rlabel via1 9 472 9 472 1 cout6
rlabel alu0 34 493 34 493 1 6_zn_2
rlabel alu1 57 453 57 453 1 6_co
rlabel alu0 57 472 57 472 1 6_zn
rlabel via1 81 485 81 485 1 tb6
rlabel alu0 90 464 90 464 1 6_bn
rlabel polyct1 105 465 105 465 1 A6
rlabel alu0 136 469 136 469 1 6_an
rlabel alu1 145 465 145 465 1 6_s
rlabel alu0 161 471 161 471 1 6_zn_1
rlabel alu1 161 453 161 453 1 6_c1
rlabel alu0 194 465 194 465 1 6_bn_1
rlabel alu0 220 456 220 456 1 6_an_1
rlabel alu0 267 470 267 470 1 6_an_2
rlabel alu0 273 494 273 494 1 6_bn_2
rlabel alu1 313 493 313 493 1 B6
rlabel alu1 313 525 313 525 1 B7
rlabel alu0 267 549 267 549 1 7_an_2
rlabel alu0 277 550 277 550 1 7_bn_2
rlabel alu0 224 525 224 525 1 7_zn_2
rlabel alu0 201 546 201 546 1 7_zn
rlabel alu2 177 532 177 532 1 tb7
rlabel alu0 168 554 168 554 1 7_bn
rlabel polyct1 153 553 153 553 1 A7
rlabel nmos 202 565 202 565 1 7_co
rlabel alu0 122 549 122 549 1 7_an
rlabel alu1 113 552 113 552 1 7_s
rlabel alu1 97 565 97 565 1 7_c1
rlabel alu0 97 548 97 548 1 7_zn_1
rlabel alu0 64 554 64 554 1 7_bn_1
rlabel alu0 38 562 38 562 1 7_an_1
rlabel alu1 9 553 9 553 1 sum7
rlabel alu1 249 472 249 472 1 sum6
rlabel alu2 249 406 249 406 1 cout5
rlabel alu1 338 513 338 513 2 vdd
rlabel alu1 338 577 338 577 2 vss
rlabel alu1 338 505 338 505 4 vdd
rlabel alu1 338 441 338 441 4 vss
rlabel alu1 338 369 338 369 2 vdd
rlabel alu1 338 433 338 433 2 vss
rlabel alu1 338 361 338 361 4 vdd
rlabel alu1 338 297 338 297 4 vss
rlabel alu1 338 225 338 225 2 vdd
rlabel alu1 338 289 338 289 2 vss
rlabel alu1 338 217 338 217 4 vdd
rlabel alu1 338 153 338 153 4 vss
rlabel alu1 338 81 338 81 2 vdd
rlabel alu1 338 145 338 145 2 vss
rlabel alu1 338 73 338 73 4 vdd
rlabel alu1 338 9 338 9 4 vss
rlabel alu1 354 37 354 37 1 and0
rlabel alu1 354 121 354 121 1 and1
rlabel alu1 354 180 354 180 1 and2
rlabel alu1 354 264 354 264 1 and3
rlabel alu1 354 324 354 324 1 and4
rlabel alu1 354 408 354 408 1 and5
rlabel alu1 354 468 354 468 1 and6
rlabel alu1 354 553 354 553 1 and7
rlabel alu0 346 40 346 40 1 zn_3
rlabel alu0 331 133 331 133 1 1_zn_3
rlabel alu0 333 201 333 201 1 2_zn_3
rlabel alu0 346 265 346 265 1 3_zn_3
rlabel alu0 333 345 333 345 1 4_zn_3
rlabel alu0 330 421 330 421 1 5_zn_3
rlabel alu0 333 489 333 489 1 6_zn_3
rlabel alu0 330 565 330 565 1 7_zn_3
rlabel alu1 378 9 378 9 4 vss
rlabel alu1 378 73 378 73 4 vdd
rlabel alu1 378 145 378 145 2 vss
rlabel alu1 378 81 378 81 2 vdd
rlabel alu1 378 153 378 153 4 vss
rlabel alu1 378 217 378 217 4 vdd
rlabel alu1 378 289 378 289 2 vss
rlabel alu1 378 225 378 225 2 vdd
rlabel alu1 378 297 378 297 4 vss
rlabel alu1 378 361 378 361 4 vdd
rlabel alu1 378 433 378 433 2 vss
rlabel alu1 378 369 378 369 2 vdd
rlabel alu1 378 441 378 441 4 vss
rlabel alu1 378 505 378 505 4 vdd
rlabel alu1 378 577 378 577 2 vss
rlabel alu1 378 513 378 513 2 vdd
rlabel alu0 370 61 370 61 1 zn_4
rlabel via1 394 44 394 44 1 or0
rlabel alu1 395 109 395 109 1 or1
rlabel alu0 370 93 370 93 1 1_zn_4
rlabel alu1 394 186 394 186 1 or2
rlabel alu0 371 205 371 205 1 2_zn_4
rlabel alu1 394 255 394 255 1 or3
rlabel alu0 370 237 370 237 1 3_zn_4
rlabel via1 394 332 394 332 1 or4
rlabel alu0 370 349 370 349 1 4_zn_4
rlabel alu1 394 400 394 400 1 or5
rlabel alu0 370 381 370 381 1 5_zn_4
rlabel alu0 370 493 370 493 1 6_zn_4
rlabel alu1 394 471 394 471 1 or6
rlabel alu0 370 525 370 525 1 7_zn_4
rlabel alu1 394 545 394 545 1 or7
rlabel alu1 430 513 430 513 8 vdd
rlabel alu1 430 577 430 577 8 vss
rlabel alu1 430 505 430 505 6 vdd
rlabel alu1 430 441 430 441 6 vss
rlabel alu1 430 369 430 369 8 vdd
rlabel alu1 430 433 430 433 8 vss
rlabel alu1 430 361 430 361 6 vdd
rlabel alu1 430 297 430 297 6 vss
rlabel alu1 430 225 430 225 8 vdd
rlabel alu1 430 289 430 289 8 vss
rlabel alu1 430 217 430 217 6 vdd
rlabel alu1 430 153 430 153 6 vss
rlabel alu1 430 81 430 81 8 vdd
rlabel alu1 430 145 430 145 8 vss
rlabel alu1 430 73 430 73 6 vdd
rlabel alu1 430 9 430 9 6 vss
rlabel alu1 458 552 458 552 1 xor7
rlabel alu1 458 469 458 469 1 xor6
rlabel alu1 458 405 458 405 1 xor5
rlabel alu1 458 325 458 325 1 xor4
rlabel alu1 458 261 458 261 1 xor3
rlabel alu1 458 180 458 180 1 xor2
rlabel alu1 458 117 458 117 1 xor1
rlabel alu1 458 37 458 37 1 xor0
rlabel alu0 434 37 434 37 1 bn_3
rlabel alu0 449 38 449 38 1 an_3
rlabel alu0 437 117 437 117 1 1_bn_3
rlabel alu0 449 116 449 116 1 1_an_3
rlabel alu0 435 181 435 181 1 2_bn_3
rlabel alu0 449 182 449 182 1 2_an_3
rlabel alu0 435 261 435 261 1 3_bn_3
rlabel alu0 449 260 449 260 1 3_an_3
rlabel alu0 435 325 435 325 1 4_bn_3
rlabel alu0 449 326 449 326 1 4_an_3
rlabel alu0 436 405 436 405 1 5_bn_3
rlabel alu0 449 404 449 404 1 5_an_3
rlabel alu0 436 469 436 469 1 6_bn_3
rlabel alu0 449 470 449 470 1 6_an_3
rlabel alu0 435 549 435 549 1 7_bn_3
rlabel alu0 449 548 449 548 1 7_an_3
rlabel alu1 494 73 494 73 4 vdd
rlabel alu1 494 9 494 9 4 vss
rlabel alu1 558 73 558 73 4 vdd
rlabel alu1 558 9 558 9 4 vss
rlabel alu1 622 73 622 73 4 vdd
rlabel alu1 622 9 622 9 4 vss
rlabel via1 595 62 595 62 1 select1
rlabel alu1 650 37 650 37 1 ALU_OUT0
rlabel alu1 586 37 586 37 1 m1_0
rlabel alu1 522 34 522 34 1 m0_0
rlabel alu1 494 145 494 145 2 vss
rlabel alu1 494 81 494 81 2 vdd
rlabel alu1 558 81 558 81 2 vdd
rlabel alu1 558 145 558 145 2 vss
rlabel alu1 622 145 622 145 2 vss
rlabel alu1 622 81 622 81 2 vdd
rlabel alu1 522 122 522 122 1 m0_1
rlabel alu1 586 120 586 120 1 m1_1
rlabel alu1 594 92 594 92 1 select1
rlabel alu1 650 117 650 117 1 ALU_OUT1
rlabel alu1 494 153 494 153 4 vss
rlabel alu1 494 217 494 217 4 vdd
rlabel alu1 558 217 558 217 4 vdd
rlabel alu1 558 153 558 153 4 vss
rlabel alu1 622 153 622 153 4 vss
rlabel alu1 622 217 622 217 4 vdd
rlabel via1 595 206 595 206 1 select1
rlabel alu1 650 187 650 187 1 ALU_OUT2
rlabel alu1 586 185 586 185 1 m1_2
rlabel alu1 521 184 521 184 1 m0_2
rlabel alu1 494 289 494 289 2 vss
rlabel alu1 494 225 494 225 2 vdd
rlabel alu1 558 225 558 225 2 vdd
rlabel alu1 558 289 558 289 2 vss
rlabel alu1 622 289 622 289 2 vss
rlabel alu1 622 225 622 225 2 vdd
rlabel alu1 522 265 522 265 1 m0_3
rlabel alu1 586 264 586 264 1 m1_3
rlabel alu1 594 235 594 235 1 select1
rlabel alu1 650 262 650 262 1 ALU_OUT3
rlabel alu1 622 361 622 361 4 vdd
rlabel alu1 622 297 622 297 4 vss
rlabel alu1 558 297 558 297 4 vss
rlabel alu1 558 361 558 361 4 vdd
rlabel alu1 494 361 494 361 4 vdd
rlabel alu1 494 297 494 297 4 vss
rlabel alu1 594 350 594 350 1 select1
rlabel alu1 650 329 650 329 1 ALU_OUT4
rlabel alu1 586 330 586 330 1 m1_4
rlabel alu1 522 329 522 329 1 m0_4
rlabel alu1 494 433 494 433 2 vss
rlabel alu1 494 369 494 369 2 vdd
rlabel alu1 558 369 558 369 2 vdd
rlabel alu1 558 433 558 433 2 vss
rlabel alu1 622 433 622 433 2 vss
rlabel alu1 622 369 622 369 2 vdd
rlabel alu1 650 409 650 409 1 ALU_OUT5
rlabel alu1 595 379 595 379 1 select1
rlabel alu1 586 406 586 406 1 m1_5
rlabel alu1 521 407 521 407 1 m0_5
rlabel alu1 494 441 494 441 4 vss
rlabel alu1 494 505 494 505 4 vdd
rlabel alu1 558 505 558 505 4 vdd
rlabel alu1 558 441 558 441 4 vss
rlabel alu1 622 441 622 441 4 vss
rlabel alu1 622 505 622 505 4 vdd
rlabel alu1 594 494 594 494 1 select1
rlabel alu1 650 475 650 475 1 ALU_OUT6
rlabel alu1 494 577 494 577 2 vss
rlabel alu1 494 513 494 513 2 vdd
rlabel alu1 558 513 558 513 2 vdd
rlabel alu1 558 577 558 577 2 vss
rlabel alu1 622 577 622 577 2 vss
rlabel alu1 622 513 622 513 2 vdd
rlabel alu1 594 524 594 524 1 select1
rlabel alu1 650 549 650 549 1 ALU_OUT7
rlabel via2 466 62 466 62 1 select0
rlabel via2 466 92 466 92 1 select0
rlabel via2 466 206 466 206 1 select0
rlabel via2 466 236 466 236 1 select0
rlabel via2 466 350 466 350 1 select0
rlabel via2 466 380 466 380 1 select0
rlabel via2 466 494 466 494 1 select0
rlabel via2 467 524 467 524 1 select0
rlabel alu1 249 545 249 545 1 COUT
<< end >>
